`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YWwSN+9l5ahBqN8tuQHA+pe+2Q7Fh9//dR3H5K2w3KRc2pla5S5ifvTi8Ak4V+dzPFwrZE+Uv4ZM
WqK4mWAaDw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WcjiphsvP4YifX33L+r4vrauIXRkGno8B+olsJNjoqAxagaZzNDAFnvGiJsIWLTLoEkntxsgRnIo
WVce53gFCvnJJkmdaYhg6W308/4ThcXkZ2dT7Q+TUTpvKAEe2vDwO0foHspYl4iLWX2KqDyY9jge
moxvN6KH420mg96l6zY=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wvng0RPku5m5MHpJv9WwJDWJ8F5PUKDSPU7V99zR5erdP7PcyDhypTKxqOMHkizg+gEusr/QYxdH
b3OK1yRKUZ44xzg4dZxpsvitjqx51I8wGaS5oiuyKX8hGtgTVrbfoHo6u9pcLQZn9XK2J/iSrjf5
dyOg2xTIXw233HzwIrCKg5RT8dfxa+iICMhoGVZIGJ68DJPwrJbT6Swg5gWMje7MS+Ppwgv0Jxqb
7HSKZuEIyqOKVjWI9mOWG9o9+LBatVHO9cQqYlFkeCwc3YeZbVHELaty1PZ3GYbJhCtr7obXWCNH
f42iQcUXnPWhD7j92uOOj9mnGCfQwEtmFpOg0A==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mnRNLVCxq+sgQJhai+B5fZRsJzZ93rdvyaCrmwTY5fIgoqSgRC5N+TQCYgevu6oU/nSzurf6krRP
lHQ0Ztrjgg2Tj4+uhFcaWXWp3gef6Qsz8XcVJ4aB4xMaBhgkUeweDC7vzOKD05WXxyBd0/qZdLtt
lS8j7xW/2WXeJFqpGaMZ30TpyNYKEPbTG0s7zfxCOI79Vadm9yVGLdGkntvGV8guzxeaRo2Qkmsm
e1+jXsDbdOr2euBE7JiOnNqartejTWUhtjRbkQnS4YCtUcNrW9+ObOoPjivEDKhArV2d5T5dFhZd
vZIU/RR6j3BExhd071LKzolsdnCqR62C9tEZ5A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
E6549NUXinEnqZcngO+xA/zs1xe2Bus1VEuxweH9iD+10PgNtRJtsG9EF7ZdZas4DjOhgJh7DHf8
ndbSlKTeJx/4QdIH6iyjSx9xrJbjCC8TeQlSsBzTcSKNDMh3HuElLUknuM+x5+UC+hkdrw0waGjh
tjj70YkP+K8Te1Nhfp5PHo+OirttOLZY7Bnhq7x3KDxVSyWnLuCBlLcRqRosb6oaQVAF5dnEKVG3
DDqNFX/V0KONWbfs5QSo5gM8f237iV+nwxPmst+L5casdH0vfnMagphcYI2Gs12f9zJ/qipttgTQ
46Pj/rGC5IRv5Z5f3c9wnJBWRVPQ0uHojBicwg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ogp/UkagRFxN6D0Tvatf3PJ+RNRc6aGWLVAuekDtCdp1urxgWDpgdUpLAqv4gVFTloxR/WYTIPAy
tqnoQwfvxF8+1H1sANWUqIMweNpcUZzEYS0M2VRPa5yH9GDRSd+LmMbbrq6RbwvXiR0tPlJ+qF//
xXzjGxQQlbn5MtTPwO8=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WS3NnUM3tGvHLrK1+gyTpPfI4oWwTOYDJPYfQBcc9ol/GaO7Z5AyMRqRkk+WEY00WrbCfviFYMzU
pGl2IHT4VRRzqqLR91kr2OFbN6OGXGirK/a2SoQqoRH7NbdhMzwc2r2DD8mzssXGs2HnjNYorDiE
Vs1axIRZ0Xwgll0Xql9UnW3+H+bZdCSjNWd63t2LxcoNPpatkn50Aa0uZrOTFNGicGTTryERIIjE
tD/W23CkHq3rM2LwJimtfOkZfT6H17TZIlmdf4GzYYEZqzxs/jkYFtiD89KMP+/WhCVPGWSzHT/R
ZumbUYGnUPG9wSLIU2c4b/c9CXNngT5yj0uIjA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
3rmBueQ4x34R5H+u7XR4wQt54c9NM54EMkf0xwo1wMnWJ8CpmxdJdf4Kg5yIyTli+//mqu/Ua0t4
++ZuiVRnxrhjhhkpHTZiE11Aj6ZHOOSrBQRDvFkLirMWL0UmYovN6S4oVQOzqI918cTMI1+A+a6k
jFweciTJtx01aJJGiT/eP6MLQJC9bQq6SGwOg+flKtr1GkTg5V3FrQUpkq/1UMHxM4ngNeYPRje1
IG1/a9BgajgWfZ5iOWEILoV2iFAWtZS8pb51YiWB/HCs50s0AQ5fKEZRt3sbbIt8buID7b2r/WTF
8FNb2xOFtNwC5UsHZ3wItlzhvChEMeqZVRK2g0nY5FPRD4lYZPNTmQRdkFPSpNWZjMV9Y44uL8pF
8WgFl4lzVj8l6lRZWaZy7dkC8TyEs1V+ooAu2G5T4TS3h0PsreLXbrogWQNw8p3kziw9y3zo+I20
cOVkLS0ojRyNJ1w/YeddGJ3pKXhz6pkTT1iAmuA6zGg1wSqZj2V2ApkgaQYIlCwEW6sWDqeztsrk
Fx3Zo75rvVieH18L0uwWmuPfebmlypn4UnNDwn5aY/dlSrxoWhwmmba2WV/QvZ58Te0yZLwE+lhi
hIvGuhFx00/ZnXE6HIoIs/4vgw/LS9zzM57oPn8JRY7w6XAU99E45ai7r8oRK5Z32vqIh0eSmaJh
rTkvg05NN4LOhf3uueJHXZLJldsMvpCc/zVBgFFzXwz8Ex54MZEkHrZnrsckK5SwO2c1T1pAmGRY
BzIqEOqCny/OWCbRHflhLetk3PkCjSP8ONSmdG+TkZQqS8/rPA7fyHFVKuo2+qdArRRMMRUg9q+R
MMqgBusrw/ab5PLnR05lnb62n1lj/FMUOBU6VWdy7fcp18PIQzH/wxH1J08xYFUWAGoFB1Ubnfxt
vgFUsE0hQ9yyBIIqUpi42WrXujHFIANgVtjGbu/zYXQPt2St62pG2AZ/Nji/5PhGJpyQSOM13ubD
OqB/pzlBmOflhPIQw0+oZrtg3wfa5bcvUIhqWWrqgLDjZO5xU3g4ECgDGSJaTgaRWyHUGnj0AMjJ
D8cbJ+N5klblBYMWCvdRi/+ztHRcl90pH51INRfit66DdEL+x6+NiU86wCSkLg5taVCUvkCKSZS/
YA6uxJ0cL8OZXI8BKJ+WBE84hjszp428Prm0VZfr0uhPvRdqbO3fbt6vxOpMelhCDWzs+RaOJnMg
ivsP1ix/gcvQHZFU5rqujbOLq0+Wk/Up1DB6YGgNcUTd4h6/jo7dhpxRnNpUWY3p4XCCfQHWiodj
8+SYnCYEpAeZFIeieDCULNstzUPjv1bigeu3d+KpEquH6i38JzG3vpc9IFfxqMbz/syuheBdw0YN
FzlRIHu04QFJtWXiTEqhAIx9XZmztRj3NZqQwtlvxvJ1iQ/ox+sEE++6tKXu46q61eSp9ARScxVa
/plke56IDuxfu7MYAXShv9FqbTZZDI0Ob3vNc2r0qAWZTKQ1VUh/MrwibpbC8Iquz0V6ttN8SS7z
oTRTxUKCU/VqOBBXyZBaqNsN5jBDs79ZN789Zuww03dYY9WunfBCBNuQGcYEgtO8V30PojAiiSIG
0n+kPWyV/y78yZBe0isOnzkdgPKXhGlcBo+4oED9AYKyFjoafH6Ww711Pb2gaQhsCgjtoR9HbW1z
32JHCCkVwt7k81saiT86/p9zGeVZk0dhdhOujlMd1UM98Mjeu4RXkrxzsj0nn0yy64Pfx1Atlgc/
Db25Mfaesy86O0rk7OW1YbUylTC9ey74WnBu2ZDN6fP46k39TViGGsQ85dbXCOsDYHBE831m6Ob8
2j7zYYS3LrhKLNeLwasrPJIZWLiL1+Q27ulwaz8N244eaXrT4p1gKFQ+cwvude4VvWEeHWJKzxvG
qRZoXd3HORRov7RuCb6iZ0xXcrYAEe6CUDibqBh/o3BzTfp/k/Kas0f+OI3kDnMrUzxn3pN08din
5EKqX6vDQtXfoZ8Y3sGNez5wfE0wcQkdL6cpH5+Zu6r7qLEuWGNp5JMLKloUYgdon0RXMJ82amXH
XkKAt0GnAs0RVcz+Tbsp5CLvVR2AE6z2sI28u/rk98UjoK0wnFtVuZW3VP+b3Y2oqCGX7RpWA3G1
z/6roP2T51RzBu1/okodUap0EaQ6QFnCw0ziakYDLn5C7zrUEKKmbWnSgvrsMK/48LuRA83nifFo
PxOGGPRFIc/oc7AFAwFwnAgDFOsoeKvn1+x0BUizOFtkrb11Sn8kNFIGHTAkbhiwuXrsb8od07+N
0CsAvveDPlrMVW9e0moW9sjn/yULgWhmhriaWTYcpCF7ckgGhbKuZx1eIHGTyVZqlv3T2cp0ZZn5
643xGjPxxTNfZhtOWkiTy6v/xCgTcJLCDX8TAgMYvGxyPT3Ueg3Ubemj2O0/5hJvq9vCob4TRa7h
srjJjEVz31b8x5yyAdNrv/WG/VhMhVG+NITEmFc6QC0xluFwbH1Jnl2Kj67d4P0fZl8TIO7M5G9i
BA+sWQk/He9+QMI1IIo6LNjBnFAPNySVrA/xOjlgZMqElYzDsINOlq5N9nxT6XptPfQ/dzt2KSCe
1FFkeRn3MNYojIOSwSBthdrFnRNI9AuGQ3pFOsprYRiOImk3HuMqeySV6xSRELvmaxGUxcaYsNtF
pgr5/Ml5xZoYbLtWdTvBuGc3Fy6p1TPsTEizZLhJYsOTKUQ4weJSLjfhpLommziSSAxbJ22iGlX7
u/JWRBheY0HwMAEh1xzcp4i/EUVshCH51FuZK32rTMNxSAl88dvEdkyA7Ea6HXpJTJ7C362l1rJs
kiETC5pFWliYY4a4iOlfO/5vfZrIYfc9TJPTBykYxefPVBDwQuRjJNHcMpirJZ86QiwI9NFfGWWE
ITe6qlDX/EIBE6CEQDlC+fYglU1NnUjwYGlpD38h/fzuzn3jQLkJn+aK0Ju8erJYx17mh+24GpZI
ZAGmkrOWhgdqs8K9soRUoBImleLbvvLUAjKsefHrsFnFcTm8uxVIPVe4RwkaKrdmHhSAwROwaQtk
OvZ68o0zF7eUnb44Mrtlxtrw6VEsIF91dNZ6DbardFqVv44Y4dj38nUhB3xb7wpTsd+RnIGJyxce
+O58V63f8dh6C3aKyUKTHS4CPuVJyQP/EohVU90+oAZ/UWaP1vT0eoJOa9S/9IOM7kKHdWgu0tj5
s3nPx6we1M9UaxPrXNKWXTn2DKvUKFbEODY222pTbUKNufkDwCYbglLqfHyA93d1Jrj7WnU6stuV
O6cn+wCyMINHDYB3rt+qHJoZDhFvKYDCXbDuH+BKT/LdAgXxcPvJIVe18osDdZPaStj/aSXXynt8
OqfdV3Sn3eb7rahaPXgWOP4dijqpOLnui1JvyUZqVvnrVwfAIcTdP/p0IoTUGBrGVPH7VDkGyh4W
iahXDWZcXLqTBd0dzqE8pV38xj3Hh8pFZaDA45MG+C+Wvwj+aoDE5xbIZYzWfhNLwIzQ6eUTiaQv
ficiMy86BhicW4r2G7FFwpZ0P6setJu6RRa2khB6d686Iq6lG8MEYlcYgSH8XRC9cz8Pdp/PTptN
cyAvN0yEirvoLKl4K8pW729soSafoK5JeRx+KKEWxKc0r6ED14FQ6/baHqB5z0tHzJfJHHfz7lJA
VSEx7cOrNRh2kToRhNzZxrtdHMFZFA67JCVbS4QkXiv+t/7is5uHeV3USMbpfe04QTmiLDUoOxT3
DwYVJC+M1qipHblGIsvxmpvZrQSjXAS21ZJQosQJLZJBkcIGKz2sagGKMj9l6cu+MWERTgdUyl6x
WMnq28ST6vr61XmArGYcwmnPJwEs0g7EdWsjFv+0X+Os/CjHPPipZowYCOzeEKjuQMPCNSk7zfZe
rFRnwnVtx1xB2kwZ54Ip4SDJ2URq2grn/aBuqMp8Hl4uWcUWEZ8zFB4uXj0A+KHpCpvO4rodiGzF
SJOCaaaZ3ZIjLPYhRN+5cF971Yly/mecFb5cuEaU1FFhenfn76EHD117JgSqpfmijZ/O5c/QccJ/
7RaeBv9X7pJtB9GChr8f+PFYLfwkcRzu8Ns8DvWR0LJ1vzG3uCSuBBdpx5R3frl1JrqL5hIUruki
LwLDfkkAeZ1D/Cx+yKUH6NN2C4J4YY9hjEpFC13a6E3uM4cLR9nv0ibFWVuqbQGW+tfgTnRDhfiw
eEZ/go/Um+QmFbENRDfWOSiTfz3Oif0hjNqW9bo/L+w+6RXo38ZR5eFMS+zK7mKmh6csakh0jsei
/K/qRVvuiRzuK2eLFulotcu4vXbjgmy1LsHz39JQ+1WoPbq+mIabSd/uvtriecaqh58CprqhU0vf
VefpZla1rsEmCw4//3m7xXUO20Tno73Vpa+Ft8cRfcSzD8PWqTPsVCrs4JnybCKlNTFJi/W4KO5g
DBaq2YeM8nz97KXAQULW/waQAxP9+apHhPOH/4XabAC/QbT0fg8vOVM7C0Mi/AHGNFztRLZfovEC
lrn2JaTPvohTcfl5mu1qKe/ij+k5MnsKNwWvvqULQTxcE6yOWdRZo3S31bRQuziMR/c6v3xP+OAa
RIC4sogJ1jag6/4rqSfk93MtAAAc0uRaICa4N3FYulTDk1oMoJ43oecIJH5942rGUEKRuvyvC7Mj
U215Sbg3DMtppiUym74EYZx5Nb87PhRm80cYyRNi/EAiZ69yy4J6mlc0idaXRl/JvATiE0TaOG0c
h0c667Qppopj9poiBRR+obsjL46uS30Za2xNhj3g2zEvwxuLmhZe4OTykr/rxUzzjYzQ+QaZ66ow
+doPmg5K7Sejch+8w9nsSdL3O1uONMLRLPzLhbiFuIOERp6y36lh+FSjAZucWlre2MEE7t35ohW8
ge+dO8VFSG00iRPllPzWXNHd31QX7PjJ10PiUAgNFXljs1TXu3Fx+LtBaHOUObC+u+tDTP3BobGu
k5FN0gQDcx2UHhrk/t+f+h0fXzmtMWvitH4OH61Hjrsy0WMJXnDxgSjnNwdneQvH9NCLafennmV4
EAEocRjMndg+WBE1SA0UjkftG3RaW77SEQVBCHkTbrWaFGHylXMvzTH92mnVHR/XwVm4IeplKqkq
l7HFxZw6CMpB3fL5niIenQx7ze64v0HdRYBM6BY+2vf9NGja7opb5qTEWiCX2It8DsUfhxM5es7z
y5XTzCj1k2wJ3mW1MHdoN1/VBGM0QSjy8pp6QAGNBaA8rENmFwAFrDx6p2WyE8L+frRemeuvm6xE
bERoN+tXtak2wPqZlfXzjcpa9tKSz52SbtWaNismbmUe6uGFViSmiwOvac4XwtOAVlj/ZFM7lk/J
gLRf+qSegrX+emRR6COmBlEmdsEsVeo+uHeU6mSEVkysH1acG/MkylU/u27LFBZEx6DijycFThbv
jHp2OEXKmcvNO3ZajDZINEglmxRx4x+r3DpW3ebpoVmgsCexbvNuAMbkhp3QOF5nODAICLrox3d1
JWf3wXWYa5RewDsT5JIDozlk2qx3fZMnyfzsWB6JYNegcHYQ5lN0RwJVrfEi1Jxq4zEu7LAcFVHF
Yul65F2ow7VXU268yRoBo5/r6tAJdNTH39ZSaJ+oma7UPimwUsH75jhC5oNShPsc4QkGBNP6fo9g
Vn3n3jbXSkd4YpW0JWeBeqTl5jmRJqL+qLa+ndG5TtVmda0Mc10Jk5AfxLi4UX/mTH+JDGDpfAAk
F8skz7B9SQdQ48vDgti0QfsUIi5fzg6fN8RRZSquefTiWrxjpDcU0IPQ3tf5zKVGUdxT0Cw40ySJ
PtNnVdLJ12dz/TDt/HgZUl9/6sFSXWITRUm1ZkUGSt4zcC4Nl9XhFQuN6Ohx87gPanaVvlteG789
T9B70qVwywcRKW27b6n70+A1UUY0TBUPDFZd/mJ9vlBRVCi9cnUq0ImxbeD6fVjkBo4ZlsnSMaM6
Ok2MPwoVu4x7Av4cvBEVrkNOc4FBb8x/AJ7b8tPvTpq9L0kT/4K4UEH6O7xWSnyaG2KDYRIKRjuu
G+4bCuDMhhVTO1lRcc0OubCF9efff1HidWtPh9+KBWMnoOSTsZpQE6gjtQeJDIlWj+uagim200JJ
a2Nmvnw5Grab4L6p5fp/dGLMRd1QchLiTBPjd5A0Ha2Min+e/fd2Q64DMfHFp7/3qprqVpZ4cRwa
RmEUsqJYmXGvIpr+kyRCCxYP0rRJ8SkPLSwFO59Fg8FaUQqLChJrUF93fsaNmB4Q/rPT65AlBSDi
KSGd1y3OTzgW6+dhzNQMpi0YQ+CZKRaGkbPCKZPs8eQ55OByisN0dNGmobZ2adU1Msm0j11OnmoY
FECJJoH2eqQFWPzQPGwVUw3ZIvAbpqMT7cwAnYrAiMxtpgLC980/H0pRmC2SJtTv7j8Stt4dMLEg
jLPF+HecBUflMnaeo7k2u6EjkkbTGw1DpCX3uuHD7rHORl1LoY7BCy54dyxVfoJjnvUgfETtZ8Sw
ZamXuvXLLp9vB9LErL5y9EOnAhXBNBT1XeXM/vjBu6FWGg1DkktMnvmgu37BNOHlsATQwmlpL+R0
KYJdmL9biMTTRdUaGPo3AZnK/s1NnrueK0InCxM8LUdFMbjqHCAkpcH/Mz+7PGZmfJnife5q0Deh
Grm5gAX2x2g6ch0PTi4ThtgD2hky09moIKaoAvVO97gSgHsglGyCmvWbb8LOc6v1ePSy8siPGEYB
ZbzKd8nMHC5cI8HCMN26NV3JmgpSaCE17Mkx14cQTMoKXlRyzrnTurwEv5STbq9GUufheWSmCD9m
tvVWSNDepqzgef0GDetn6d5XRBPl+R/tu/gq8aTb6TaGReqBElEIIFLVo8ohVEduk6tmd5Tbnb95
yv0K9maO58z3qthQt0PSBKJ33aNgAwktkSVVcwU/t447DJwhnzFYFGBuVmztEGmyqU+vy9wPA83X
fSffYX0v2F//4rmXgGHp3z07Umqb8llGx5GXQ7g/ihPz5fFnXrsgdJHDFSrEFgblmGWhHfElAGNS
ddit3cf5pHKMGKsdOP1RbPDmv4qFIKH/leMEY95cZEH32KDfqGVD4PPf3WOBHPHzkhkweimbcojL
gtbCXXFLIC/lALiy8bL20YyNdJkq+1hP/Qtm6Hw3t1u7tuC/7q+xHKTw16z7gXwvgkWY2HaSTWKo
4M0uolArIp+Ba2tvl7aKLYZC64uuCLsFn/VT4Ojqb8Q6K8uGhWnOD09csc/4bpyvqoCfJE40ncpI
0l8LSaGu9f3HV68HrN2dqHTu01QddoIHD1lXpbyNIusebW8g14HB9lrBd+PakwxbyINjbLLpYoNa
oOVEH0zfAKL0spNsICeLsV/m13Wph7zSsfwt6iFrCVwthtOml6ki699abXn631pzYff3zikapFxv
iABFhQD9V8ddi/55Rs7vi4S9U7kuZd3XD+DTS6jHwBeJL8IbA6udii3a4XUm6XY+NTNK/9Y2sEV8
8DyHBGPG9eyS4tnQ94d0qd5vkl3nnpCL7UWYC16WMOLSfzbUBSQlqIkUcF1qBhQ6SVlqP9cve253
/hOrq/ghMmJl50qMMWyNwg01WJ2J7/vgZ6hh4mnMVr+Mn6AfC/unvzauXishsJKLolFuTHn2Tn0p
vryMmJHEIQJ0ZxK3Pu2Tt+zPUIfKoMNJZIjpVghI8ZAWik1Lld7MkYS+FbxSUWVU2bJxq4FrvFZq
69UCFLUKKXFbZxJu98X6E4CwMvrBQb9917VReIQN+YmS3PRep0qkognEkXK0Agl1mgD+CMdZgW1x
ftgn0YgGqRjr4StjmKwvtOduogeU3mfR6vWngPfaZg9XTqsEGrSJmaBpH6Howx+0UGsl8wehn8M0
3WcW6CO9NCI7Mn3SjXRGKWiI14ONXBjVnbHz2kIgdKYmDkz1yKrH6raz8FOxrUCo+O8e796Si2uQ
eBb1VmfnDzmKe8Ug9/zabK8y0Bob2dqCGuA08v/Q+/W3Rwb/DAx0DMapzS1nynDye1uddi87k8Pd
460Id3RjHPcyuBt6isC2+/eE7QWZ2Pnq4Ec3PulOVT9xO0ZRc2vHCs0SeI3FI3PsDZAKCpWG2Uuu
MRIjXTH2wMzmcsQ3EKzAQG8+Ys49+5sCejyxmRT5IfCz77jXxSoFYPChKckH+yzKIMwtzMpsIMg7
nZ6tcEaCEsRswtM/WuQ+hz0sjEVdx3tztP7XApWYFPW7vA/N6A89nyE0xJCMhBXS1NcMIIswLKGn
y0GFLHvOX86NcTwTxcJWJsUmM7gv+YktuzSDSVcY2Uiuf0KuYbz//bLCuQpNbivg9BWX/6V94IX9
3cjnAkGHY3oyL1wLAwl8qLp++5Hlp49Iv8/L9leYGZWBbN1SrG0YaejNwsHv1rvJXDRVAIJ+e6em
Y7RMA0D21GZ3S+HuheNafU0QjrsX4ib75izk9niL2ZXUqW15PV+fpvzvTdwW50kNTsGnto3tGEPD
u3v2U29CI6nVKawQw/rHr3bFzAMrVHSeanrvimNTWyCN/O5MO+gyesEqq+lYqtGYJlaP9ZpaEAyl
oVI/PfqAX9TZni/qEPXrhE47WUg+MYWO/5WShwk5OXCmEJhsC5DXKG26fNR79hyzNuNEoRlrP9n+
v0KFRLrTCWW04us5ys2N3ReubcjMUOoiQ7ld3qgnUgEwLH7Wsi2LKlxUBmEH+jKEQuIvhfffP82j
EOGS+dw8+x7m1j580GxKr3HQ74uQGsl6UkxkJ8AvY7WObfkQLWmEdf+oh4oKXfhkhrRbCbwhV6gm
LwiMOQ235V/Ij1Igr62rqJrNsiVQU72XgMHhKqGNtBvTYFl99wHBaDlFjUO7+CIe3bRidoCDI97H
GnIYydoyOXwGkKh3ru1QVgcfLi+j4TvSwrM0SqzQrwf8DbL0ab52TuaWyrE7tTU2J/C7VDJVrf++
ixFtUDngDr6epehOXbQl1ERx7ppUgUF5aSDfRtztJQBrqc+spjE/KaSJ7MQkX6xiJlgMaj3e6HTv
OS4GjxR57u8B9zcFwhKBF+UlVQIrjr1bPwcZB2vEold+ej6l41/FpkXJVF79+h5ETcwh9/u+gUck
HNh5pECHJ/j9BP7OAGoAgeKPIckPIuc78afIemdOFBaVL30cxedgsG5RIdLYfzoy+3DuFLDmkhwV
NXArOy4OyW/IJwr8gWBd+Aawt6lnhHmEoaoRawIkeTGijKJPTquNgfKjEdpwPksTUccO52IVButr
WE7Le2Ss+hmgZlfnVc2g783m+47tOGQWo/KyfZXFR6N3Q4wa+IyXpnFKkpzBZ1Aem3NXQde43u8j
8gCUxmLk/04yI5UxHbFhheMqPLO6kz1ZkwbwkrMkI2yxrnccEBFT+Hk+aihSuided10xLcd1liaX
dW2vCK6vcpSTI2pZD8oBiMN5639innzOzXEuT7RLkeFjYpqhCXboU3wQn8DzDDe0K40xS3CShMWe
Rc8pGSS0B980ee32XDkaVwS4Z8X92UjCuj1c96xE6gVeFTXuMuuyh43llZcJ6598xafier1NR0Hs
TwvNveY9jfwFBfwKVoLQLGnB6gcatC+o3fvhHDQEysHj65EJBlhysyw+u03NX2rMcgkXRMVb6VHp
NKjjlh/A79A8uMLhHsuxqR6t6t2Ji5BJrm1Vsm/IUDQQemT1Qy2Nq58wylGAfPSFY+u7KiQmbajC
oziIfkKQK+oE/CDDQhZWP5ns5qIIjnwD/4BS0jQlvo28+V2LgplGyI27WxvKsJoYHO2qKKFzavgG
LTQcvI3LvWwn1a+vQ8IcyGKlgw3IgOFAy5+U7fZfggE3rXGVObvUYU2UuTaYz1f/jzMXRqRV1nDB
sJ5aVz1MAuduWpIKVigdnzVTky4x1nwF+NKVEkDkReLe45cQvr8MXiP3MeGX1OpkzBVhQooVNPSo
RTYIFO4SjPUdvmFlwmSi3TgDs+tTD3NMyZILcW+VqZ/2aI0I82dqaAuBL7j4BkGBKSI8Fc3FqEGK
7U0zBM+KpXwChqNfFNIt1wjlhc1J9fuDcBKyu3rnpQPMAbcqqFEMzQZwH42XopLl3Mvdp2i3gyTk
9+kueMiPuaKGOSWzMYRoBLPFqeDI7I29r/by2+SHBr29bJSOhbJpGUrL/onA5sOWDAprFa+XfE06
SpK7nxmXD+LyJuVX03P8kZt2l/Us6uuvZ9zaA494s2JnYBvYs5D1hJ02Qv+N+tEWdINohvtpEBL3
L5W4ikSD5vkTSIdqKk0AYWSJ5PvgTKMrIqUAbQmKMYVLkimgY64+kL3EkzsUi3GXdxYO4OKhn0ug
QuR0nGjXfpsXEJ5ZuDYW8Q7eg7C+gkkgvEb4WIs3G3V+PuWCnl07GL+x1bwyfwBT1kTVN82MUTVO
EH3D+nqLXqLOesJ9Axd1Q9eEiB65TmZb/8OFqEpSKYJINIzIFbheIRWdUSqWvlqzUCKCkx3ZIL0P
kQACadaOpodK44pUhIL73UuiogVq8aUgP1BzVzpgzKF83v0TRHbd/GUUYGSPVFLUwYRO2XQ/mk8k
SDo+79MLyJrvVbvMVLfWkhwa67JtTa3jml5HjGcH03V8McwKxOt3MsSSX02RjnoifmgDljNg5FCE
0ArU3TRC71Km5/jc7Snx/OYTRzhD7O+R7EOzCai3hoJaIHrWou4uoePjPSs0bPc3/D8fvsKmgn4G
BdO037rmtHHQPjfL+jhcblqjl675dt7sffxqRQCblhSsAIdR8KtOZLq6zc/q05Vb8jkj24h7uvK0
SwTIWZLlQRYv2Kz4qN2+1Iamn6i+azJZbvu1WaWmuDVfcNeQC4pYKs2zjrBY/AhtFBQIjxkjVnUB
Ec1GGN+/vyA4EyMMPVrQcxxLtlGtAjMyP0KGzT1tZcTkGOtAkBeq1Q4MI+Avw41rAP9Kz0d6k3J4
Vw7UVOWyCjIObn2/yVXfdJlMu2CjJspUP0gyoDXXeszFg9eiZ/ZLNDqP1jsQKGDc8xeqJr3ZzE3v
NlGjO+82Nc46EgV8ee/hgmGEzK/62tAvzpPZJ6GPqDN7Wq1raKV52vnF3cvOKMQxbEmowzLFdtXR
FYwMs5R43fjmJCgAI8McENFpEOPnsI0Tb8bT+UwFFEZtbp2R/5d7INKjCHQTqKIMcFr82pcnIk4Z
I0rnpBWjg9kfz3VXCormN5PFUdDUhHFTP8TmAvnHo2om1VVSbtbKBVh98E73cc3OR5wjHpzt0BwQ
Ob32hHZW4tIfuVfqumLAP3Xsnw1nvjHRis7O9SWxGvfBep1oEFPiF5l4hx+fAIlOB+NX3eQRfGaG
yVs6lDjd965CXoV5q1r1RdyKuBWJDynlZ/fcQxubyeB9HD+E4wP7R3sq8We2JUGEDqTIJjkBB7Qd
PHQx4gMjuyXNh5QuRxRqaXlbTFGCTGG4JNl8ZO5btSSU6FbEVdKQLhakPrZ/B7xi0EOVqf5rlqdF
IPleBvMf9+h/VFmIURVv0YjC1rnbeQ9mr+Og00nfyOFWAK4uFu6y65W4suxCshlbdtfPq4Dreucq
kKSl8qhbvJS9TLrMPlq7Tq1eFfDARU7XvR1aUApY19khubBE3xDlqDiSGO+cEddwziXHJQ6NAmWr
3JLrlAS2EuQvdRbmcr89xKHA0zvRDkDfjX/1BMNbfiq5V51j3ymUOkKYjw4ZuOaYe9OLphKo0aM/
eXTLpIj6ORghCe6/jPXPheJr0JNvYbPw52oTa6oVWmF4ScFkbrQ8qs0etP825PXH/kC97cQ6+V+B
Sjfwvq2XiUfucIWOt9lOmUOaodYZPnulI2hGtHIZ1w0RJsMNKA/pML0u5kPGXwq3XAQNd57AVUxx
c60u58rRdVLrsKhrgKzDp+fxKsNQqKlWy/PJNw1CalYE1p8LMlgKnWAfuFJEPjhCituImnuuLuyY
d2QUuCJ2yJQTWqpN0EzuFkAJ1T/m5F6Z0WSFZCSFfkO/ngDZ9A4lK52VeRLLC/h7x1KQc4o0hDgY
CIa0lkt+aWNh9cbbmTje2FdsfqV1Fy5G98afSKreCUNL4zvPoYm09rZx22If5XXRfr+bCNAn8/uu
0xKokbnb7k5ue7HPnfPUwg2jCySivcWU26nyY0K+WFNiyCcBdrfaC5gFtayOzDW+XJ62IKZ+meLY
Kz3xPUGtUzLR/o1hEzG+LaYnT0H1yqltAo4A4lFOtinTFGal79jKpNpHiYlOCbwAaTCwXKo0ltuq
JCgaBqn0L/Juw4d8kqs+osuPo8mW8Y3gjGpH6sk6NjASiDvctV6ud4L3tlsG+e0j8bDO4rDovi4L
hqGuK/kSzbtVvNt0ZUV+Ig71VudqCw4ZJQnTlo+eKqN8uyFQNJAsMpHMmINAAQXhYPs64Twn8SO/
lecm+dEINB9nKfB0P2fhIAuEYzCyyr0aQLKjQRNPvt4ORkdN5lVKiGZeNjItRn5l4rU1Sv8fOYQG
mTiL85xTmCd7zfxwP2iXoq4ROu8JXv+XeqdIqcaeBvbDqcOUZj+9w2ITlfGbLv4BKjtShcLsWPYs
mSV4rVYeK5N9ghj2cTivHYf5IuujxBsSePTPYOtX3xQhp3YAGzgkRLXgy3YSjfCXOF347hixJ3Ae
iiNTl+0txg9/azUEZOGuV5H15JYOzXFbhbUZ8aFJw2N276/QzlPV8uX7REcTIP/C7a1cWyC0HV8+
qAJ9BvJxY7KID8foLo0D4UNT1uj6tzX8s5AkE8LYy2ot7PdNCFehjkIIPiyzr78iJaOFYrxZa5U6
MCUPtEImGQ31DTFGHEL3nKiDCWSVCF0vCtV29BvdvlBNFtyggHU0a1xXxgZR5TrbAyQXbsu4gcgM
A3MnzISR5VpZgSgkQW8ruZoAxEm/BI8sT/kUe2N4FzQJvtFemMK1ahVANnyu+3tFT+NlECJRv4qI
i7faMnizXKI72AuYPx9oSyDNY3FFwKNP2HzgG8N5CldJPaLQdFYocbY2bwg7lpI0SpBDZXpzcoxa
cRjgXotU1atOs4cmMwKfOOM0kLpD6y+bx1ZfUch2iTuGZ2CFDNquetR6/VH+XBuMCrYhuZkcsKrH
+ZpV3kkTYiqHpZQIbuLkL2gT+ROjAgu+0YIQRSS+wECLPclsZbcLq2/D32CuByreUSujWTP1JxWz
e6Y8kB5eAm577vqFHtzz1JMxL7sBzehRjTdjC9zIZxVxebHZAJVnKT8ho0vXomhAa0k9l2IVMPCX
LMWIuzSsayXzKfRsg4m3v7FO29UJDRbJN4PmaQO+RPi9KG1fi26bljMCQ4P9S9SqjQZzfTKZqw/p
0l2RdD5zKTGdqyzwKGXhhKc38yLFDjQhObrVbe/qg1RdTOYMOZRT7Y/pVuGLiXFIxYLTt/Yhlu3x
rDtupGN6SfKWDI7Kv8J2kNVn5K9dM7R8yvMxDjHUKiG/WY7HnFRXIu0FMDyuOZ0QIGnOnDjlphiI
iQ9PCmgIX4sqj4gl4zWH7/5ilZThJS/WOirG/EukOBiRycgBRhRHbPMy7vJwMoOdwvmwUax3edyf
nnDz9VVG9jGG3u747CKhg77Bpm0VlSDHebM6Wrz1CC7N+Cvmw6hfzZfMcehcVR6Cy1GkKCGTa6fn
q/GVpIagmSLIasyygOeELH25B3j/ONGI1iHhB5J1ma2JU5RLdD5UBd7BpzPTq7+1RevglW/efEyz
8Bgrwb93kNw71y03YifEggBaefgR5a0EdtmpYekKMjOp7yhk17e4gE/InojTIGZv10ZZBrXBESs3
bt8q+wjqFuACcAdWtNkYeuPzSqZJVQ37gS3xy3vU/ck1pfTn/8NI2ELKZPL5J17JDef/RnHo4cWJ
XTzR63TyQLEN5eCRfH4SMnSWcUtpNBAh1E5H0IM8UW7hcnMte1Ex9MPHVkFIg8iOxuJfAaGm4ANm
o0IHJReBNMxPQ9KEr/7Xe6Ojw0qstU1eSSdmwkwCFmTV27JPYTyEcjMrDUzXnMSbejNocMgG4bxp
tSkVPzJxqZDtlnDoZBZYu33MJvYV69m90XriZAnr4zFlyXMEdRbIghwDwrQ6+K+HQcdfbrPpij0/
OwXaIW+v5/Iv2Z+tWYIu8xrdRDCLDuK2+dFh0CsHRA3WFc+GR9QYD0g0P15rQyWnL25tCY7daQA9
Z+0Yi7esSlDk+ihDaNCerFlTy9DUHHvCAsJzonfvO7NNaBmB253Sef9iRFsi4Twdn8dTAmWeaBao
0yu9axpLyCMCP2voPrXBjpPdQj/x2FfFTAuPZdVrgNP8urqHLStdAkgKWH9GdMZNlompnEFDpR74
ZtC6UHTi284GKjoXuMHxNAP81D98oQT/crt8ZkBCJm8midVQ8N0fngN9vcZi7vapq+w29PJyVATu
NMB3g8XLwhI09NaqPL+SM013xquNWsUqBdcE3HGQnlL++sr7Q01e75/o6rLmMkEz1MrGyLch6kqq
3AC39Ac9d5JoXOLBmJSL2xJIUCBwlsIwImHEmwc87jxGOM+m2pAy3WF/s3pwrWwI0Pb7lyu4+J4D
tYwQDApl74VmnNM/2oNlmMBjjoV84PW8tn9nw2JyZnULRmdjp2asrMBgoTKHhuWa8Cpu/ELUW1H8
FtkP3V6qV89oXrdIUpV9+IfqB0f62A8OPndrvXk7dS/O3zqGwWsQbtakKUlN+vYt/qIhiMapy7xK
nF54D5dW3gcfPnXGsX3LQqndSgm5Tt8GhdWpYgsm+gF1padfQtltlZPq5LL13vGm5v9rSxez0wp2
hfZt/bB7IrV4FG6rjAO19rTjeJm3J1ObbZTXb+Vxxc5B03+8zHpqkvOdl9pGhKS4hKP0a4VAa9ur
AWoGWAkBIaSYywEtf1qnpsfrOIX8poApFbLjpTKVY3x0lqmnXAjtl/03G+w/xo6jEOFmYWTGVPty
Brj8eX+iydxUUjj4oG0JVP9Blg34/SjbHtk+GosxgWT0C4Rv2t5yq4u3bJ51PUDLEjgnygSMruAh
PsYGjsAjZ6g+4OLIDr7f0R+7k58nRugkTsyJf0lnZIuF8FG10dZbE9g82tsXVOUHCsEcmdeUt9TT
NNTuqAtXZHbWI8ah1HvGcmYefJz1UvoxRUJFFubffKMDwbasFOjBe62xxSI6IIWwR5dANQKt0K3n
/KLtciGNoVr/DBgMmkpQxpemXOqsz8jqufrk3RmHBS9qhyeSvCnUzajTBkXbSejqAWKp2AGji8ET
Ne73teoMMvkVkGu9SGMkXICAQUuQTiL/9lp7h6JnX78wvnzD9k2+8azr22FIXg2sR6DSfaRkzS0k
pYr7jrsUEF0sF9OI4k3Ga6W11tTb+WoAIpKfhu26gmSca5DvBH5neakuzRLZwfXvvlrxT/qONbHn
RaLq+p+vb4J3iJNzYCZCozu3ClVbKxJ8mI7XcyFW+o9Hr38mI4qcTuYFKHTmovkAjY0iTsW1QqXW
RzphdA03JyQ6EUwz/yTm5KLrgU/fD61rHYzCvvIdkqetaHgTtlkxOKWL3ctrAgVFR+pZN09NIuBx
MPlFQt7B2TeireNvakJO8PmOvu8GvazwENReP1haQtNY1lGA+xR6lWjHbgHxoLIopzP1F8VLd/Dy
Ih2qLHVxbiBe+nBNL6gltD2G3Swt4OAsZVTTjpEfy/8DQy9P9ViOTZRYrYZ5BjHg8y7fTX/ZOFWZ
SIRP4MknasF6Jj6uTmagFPu8Y5XRztuQNxy0L8eMlJTxc3dhzHJ8qqj2J3/0Ke5fyWwAEu/Dae72
coHJenkGdNOkG+MF7nPaFuQy1W3B4AtUxOhaSYvDmNmXKPC0N8TPztI6tc/LyLpTuyA++rKPgMaQ
NGJ8XtYqTjgjbe1oOZZ9CUvMFFhCCZAMkrF5L/48MjLCmj8FrhzShe9SLNf+DdWoKfAQiU9GSfGu
wA3BLFpmyougp2pRqXl1Eijcfnh3CdOyWIML0Np/04hWzOm/CcpdRaE1JT/+21s8ol67pXphuHGj
5Yc+f2oU/HPqZqhuWQsVH/3H7crkQFc8J5kyIYMiRjrUm1OxJD7MGtGcORzH57GGJq/IdluLp/BC
Hith8+p5yialZSMj4T2ybYooC9SpD49BeOwewCUyduXWxw/JPsfrLqJpfvpKq9e0CS7pQEwRXhaP
vlCt5qfeLZTh7ju1fe8+fJmEfymxwQD83nLDn5tePsrYdwwyGOmlS0Ds85hvHyJOLcBfVcGKjCQS
tNhEki4j5PcOuuo0YfRYq/Z5RyQZ/bP8Dy1oUXdd4c1iByluxlD2o9N2UV2A7T8IwvIBseaqrE1a
gVbHGJelOQR2lXUtUXgbbTMnCdFvoLLgW1vN5rJdOEtbbPHe+B5g+ou7jAxIAv78/ylSxREdme4q
3mJ1JtNVpKf7qBj37FNCJ2j19ikIU0TNOQWjXdrGGYkpiBuevWOLWlawkuwWZQszVYenjZhG23Q+
UDanET484ldqhLimzr+6QJu8yCi2IRRptMyB67PoJhVVABr2t/XlaFRkhkCa7t3PPDaT8FbU/rUh
MNrvgqFMDD3yrUjmNwLp3dH29Hv1MzqtiD8BWos5q0TYtt2XNyZF4iZHfYYbpOoZHbo+B0C5KCMG
oqrgRiXkYHvr++uASp5ByNZ7xLR2AdzJ6TvXSAk6/npZ8p5G2Q7UdqmhoMpcq258ClNbCQDxGu2r
qQeueJi1YOG0hENoGy+J1tIvYgpdT+LepvDQZRpaL5CNf7GPSHw0veBiGIPbrRncf/1PKW5fLx7I
EFdJuRm9JXY7NL7/oZICczA9E41QcVIxaecXn0IQ56SU9AxMtvnxE7RZjTEvGaaMb9UKSzmcZfGd
DPgJMfwREfxSOFyasSFDmIraaGKAK4JLU1XEmklzl/zuN9ux3H5eTZ/xmp5SuyukUxogDgEz0/FZ
M8NGyJO1RfrjOkxBUEMQiJRY+NabbbwltFlMYFtKjs2S7TAbJgMSPsXwuRT+vNcAwt6QNoWwKxu2
9OlFf32RAwgFylJSgejRAVgIzv5o+xz8dSynDmFm8PpfRI/MQo3KaZrR/X612Dhn0XVf2/yNA+bS
87qlvb3EpgdNEgFPFMqUQXpSLaLGNCj0jsGKugz/8YJpCIGgupYPby2+H21fPIwUxc9VTU0ndfaU
p5RDtQNTD8RGDLI2Txx2VTZrTBng+bVwBMmhZOfWMCCQav3xsjIIjkCvwAiBuTu1Cl3bwy152+OI
FPX8Aii0aYOV+0o4GJ9UyHyTHbJvhtR4P2Uzdn4GUmfAi3aUzh3h0Vt/aaFQ/AL3GGtLpDBABejE
vYW1EdDs0hQQwKzyX+z1toDn8fgsJLlpAiuJxl4OIiNntmjgKFl2xCfVoMEwG8ILH98O0PS9vpwN
PskfbsSy/k2FIsIXqMZWjMIAhtasJMTtN6g6h2jp+CJAn5vj3AFw9BnjvGai/dPNjveIUk3LmmrY
UoC8dDryTZmjA7uSwm3w6Ch64RGNMGbOU4kkgV1GyspkbglMsVWJm7z9lOnqQN6LWGSBK5i6e686
EuMPEJx8Hd2wQYAc970FxUmByWGofPEXLQybLo+XphQkMOwAH2GPysod1zT3Pz7d+0jLdMCggj1A
lBLpAFR52BFvVu/y/S+LTCbRVHWspfG1FLTmqhaOtnGQcH3SeewWTOE1tT+rbC29Da9xAA7RgR53
AofEGM6MLHaqeSsqnxsslav05ef2AalX5+JCUwB6IrsgtaTAoIJADGtOJ+GyGu1I1hvaw8ytOCmH
JRZj5AeyfztEIlYSmfKdNcpwfdObpA8iGeBx1qZRdGBMsY/i2slzLRRhr1U7tAvquBRPibZNs6iq
ES9VWhqFYuyl/Wn6x45EPVInAlTEHUnpLdgfM+XzkMSDmixj2VrQCRjY5ZYj4LhFBbnczuUz4Iai
icXJd+dqcnfs3LrXqRPr8zQb/dVGCtajPujjto1LJKmJ6uCevgQ6s3J6xfYTNt0ECKArs/8mft+u
DYKQYN2xcizHM3sVP+WT2M9RPz/ZTIB05T6zx1zyV0Z+pdDp/uC6ghtLu2Iqt58WWCS1l8YDP5Dt
ohM2bied3ozXQIHEZYSbk+30NzUqUbRiH9It/jD7cnX5Nx+DqGLm6V40dddXjrQ5i776mj9OdpgA
h60qzemA7AuD+9wgn6OhjS5DQUp8e347fnX7h87AFyMUITOPlp+rhprDDmdSqYUnEF1iARC1aPsB
47DPQWkZcCtESkYS3qvlQqQ0W2dmYqluFxlbvtvCqVeGi8kaDz72qdgtuGGcWrMAiBAmSncvYGjv
OOnKGZ7U6Ohu8jd5JWAFQaiSb1h8Nbdxv+vddIpQx2fmtt95vpIXprnQ7Tm4h6/zhJK3pqzkD+OE
tg6Af5R8TnjPjHSalBRaPm/3Sp8oFCcEzzrsL+xgnFshOEDY3UgFuzyCSTpNfw5WTkU16xuRjeq8
Ztb2Bx/IoTiSedFKZwCVBPCHdGpHHTAqm0LUaQosAMZ6KZocusmT9VraVvBCtqUGFxL2CymP+PwG
NLpSEYfZDAR8w/ItU4Z8de/8RagZvVEkd815S+Cxl/wp5sdUVxNWK29iVIm4SiC+eBsQGFtbKEaE
mn3b/N9ELCeoT/ut8luJ3yAEG039ttIoDHF6IWwBr0JQr4sXXkjme6b5d5rl32jdyoPFpCS6xoEB
7G/GTYiw6bTzw9dyU35R5gUxAy5fSa8oWhJba2rU+nyj8NWfCtk1juH6Jm3yiGjUNwW9/YG61PsR
QEzvJh/Wxs2aR/gSdakxJ/NnxlasKNqCKdWw3tSKK+LmOnA5AeSvpytm95sOiEHybYUldckWBd1H
BuqjPgFsdydRbf92QsUJE5R9wrYpu4Z/2W+WyXDzboLBQYRBP5L7z6lG0ap4mfVm+6cDyjHBnRhD
V26jZ45sM5XkTyMENPDUqBAC8vZQj3yXFGQjx3OmGOshyqt7eYlKBLVmIYqyEpzM1NEjeUpX3Qo0
dvQsRBxO8FKOMtXd7tNee64mzjefJ/o2cAeBDXASDtfATj3StxOyLDhYJSTZNONlqsILGZqbjVyi
NLc+o4bubeq4vaIcmUIl/GdWbNXmsAyt/1BQ9iVlEjvqTRauRSaKCrFn2Tx1bjvHtP+aJc4OVUrt
tNnKqd5VIy4a1UsnBi6AniZ1Hg8lNcQlqfowNsgX7zNa+OkCtwllLdHhdVaghsTPOSfo65O7W9dZ
/vcoMrP3sJUTyXSjB8u50xH8kz9SMAFmeRsUNbb/8g7+9vXPMmAamlcD4N1M6l++R88dV5YKQaLr
uN/v/WG18KNyWUjzlTjAH0pi9GOYkAFUve0Gv2gz0x9bNy5gat8FvtpCRHRuHvY5Fgjqaungu9jW
COnAzjrJmfp3A+JpRWD2Gmhc9bsUbtxBZgPYH+b79sHp5di7b1QpW8h1PDrzL1e/LOzblHyJzWt1
TPTra25AxRQiW6TQihE/SMi0kmaefljSrjc5Bgu5VCtFswW5z/IKpbm71d8KVVtTU2bjyNa4s9iK
yXap7u01w/5Th/Yn+V4vfeYsNnmBnSWD+L3+h6nAJ5Vs0gjOO74/vnrFSYexFKRESCPRs+ffFvLK
dKz59xyLLocVZJnRC8ehq0n7fKMZSKKVRsKUoGTM81n6/Fm/WVyiaXi8RozqaIcnI7Mss8+xi3Ie
XvqgGnNg1ifCEBulveaqqbdn4juJnFKJfIGjqEqmwQGuRl7UmpDjQhYnVcxLRtUvVHRedzjkoH+Z
6NHRmuYauzmaqIUPixcjSESj4qNpiOo9h7vfzUzLTEA9VfF13ShDFdB2PWq7JTTEVrHcBVv9nViE
kYfL2/eBQ16ogIOwfQAB1xe1qx6h0oi4/Bsv6Za79uOceICmY8aRQ6fxsnDlxtaFPQSSRTYLv5Eh
DxjdRU0rEh6Um9VQKVUS1MCfITp0FLfSzvZ0sU9Of3LCsbkXBrcLb8lUcnuL5kPIKUXZhS1LG1iS
dcCXR309Xj2oEYD1F5FSBh1587db7214CbajA9cG+n2vE1mWxx65z2vwqbG8jUdWgVHxuSupjSJg
n2VIxYjc7ol6kwHb+FXykK51NHf5jZOf048HrIxH7PAGQOdzZ0iosAz4Dj4jKYGhQl/OASuQD0rf
G7Il3TWEqj21Yi0V8Zi5G47JdhMg0xZAX8pYgRqwBlusVE62HX9fzm2duFRoIkVHpfVstwkG7ib0
jciqetq+Nf2uE6uvgwZegrl+Frd7h9rXdBMYMZPhBr9Rp0UdfywzwWrQQ/nGciaiBUWJYxqsqAlx
5fEW7wRs/ZvlQjEWealyju0J3KQw3U3YWVXbTYErwXjgmu9++lckI3G+lJEUXT+vhdNo+xYMltac
aPVgg+d374H+9Lbz9jPzLPNzpODcE5dubWdCZsPvjBo1vwwuRMoeb0N8A/aH26FUqXAWLGjHC1jL
jXzKrkyLQN8KvfuCMZi47BoQPWkiItEsO/TM/OEB8rT13ko8tBQg8mpg7CsGB0p+urr3bICaNcdL
ssAw3oN8hh8td3Bvjrju+QChvTZ8l7LB9MtXEiZhENoegY0p0w464OPLMs8mKT3+0fObTzVoYv2m
OgJ2bxIrQcBhZNODAzZjKbSTijLAk4IeXym4YVfdxerv8FchrbqLTgR9nQ29BXMENpzjklEFEh7q
BupzebS+ekQA43HD9qBKl3hR6yHZYbUZonbjS6YN9dWecwrQqyrCoIhSc98zi/MFeJs6GSRN9VW2
9Lzx4o3rCAflrE0bAE3JZg7arXGZRCfJN2t2b7nbMAhMX9RKS3xxuV4M8nG4FwB5y+ztEcJWEwBx
1QyWryYyH8rDG2KWIeZ7r6kcu2OIqVfdujYW91gduDrHg7WYznuYFtSdiFuXwywpTofyB4vzBeGw
KmjCJE5uoHlc1aMARQ9OPoQDm1QlZ6V8QwsQdPQDpDC2MTLwyXPE7e8xQXu6XrgNTve2PGEjL+Y6
acFxE4cx8uySeQph/Q1U0Lou/jJtiTG7h6rdt7gsFmAbV8TfR0wmZCxuIcrtvln0EZZ1q6FQcc58
eDqR13TDt4jzsUNM8fW3xWXgI+ymacCfOQO4ipNNpcl2/zzZVSwUTTK2poD5qAeasFj01Y5y7PDY
pudKHXSE3pNeh6i1UkFBzVfsydXV14NjchHIeHnYo4GejSjrvhcm2ttUGC4Oh9rruF0lSA8byFWO
VAccpFmHd2Y6wemfSlBWhQTI0WZrkb++kvdTs9vZuHaqPH+qZKoRq/Kvbl015mHau/UQVWv4c0u7
c9muG8rZvJD4/PYLEmdK6RJf99vjqj4qNJpdbnrlgmTACkUgBU2SUE3Y3beHiF3dwrhxsyzqTIyM
HAy+/lKcWXlpqDfa/q7wrrItaqXryxr4+lC3O5m0Bi9W+g8j3dHpSnYsPl4dFY8sdmAh/7IgHXmN
GqWhhGKmRFTS+f0OqW+Fo+jmrZlWTzmdfphhx+kQfegbgoko0L+q6IBwlXOKt6FO4OZ/SafqYaIq
scxRoncLJO9o5elcDcEv8k32O9urkHNLLCjp0coOZJLKR82uC/kiL0PiBTd9ByMUObqNKPWH5Na2
z7ik1JH1mWaz6dAjVS3v/3LRFSyTaWVOoQKah+9AL+sg/X4QB66QMuenN75BLpna+RAPQW7TPNoZ
KgIeowHPyklWO1AQLPpjuwRpmJm/l+MTjTLyp/4O/Vm9R1HnmQ4S71Lnr6nZL9ycFIGO6ep8BahS
IZYhgqV778T9wa93E5s+3dO3Sh6xzmKKG2iounQhx3ab7/+phPdF2jLyx4SOrrrUYXRvnw0xW2XJ
2i+DtUHdE3oeLeHHOYrybkp9pbwn2RIqh0PEjznjJDvsnGwfMMZjSbZ1YGHEDswqwPeDHsNDjgfE
xCcaLLYYQ/odgem2VS4r7rGQXClYpPMEoZFy3Pa9PcXY56CFrjpNzTSmz8IGRyirtBWT8JqQaRmt
FN5sv8l+P92yhgp/ZMwhSbFB9SyqTPoVN4KAx31+CtMb6/DxjqY5zqkrRavLKvDUsMYjsKOzwwTN
e3KPS4igQDteagjGJp1JM1eACWXYba99ibOdP0nYvvpuDVW8crMefO5hdslwd2BdLLOzgWqlLrtI
UGVS30b5VGNBl1w9Jmj7W0nv5GomQCEDCnW20QA6zYyop68Zg9ML7YIWGrBUxAwLAliBDBfrnYlh
G0ItAEnrmUZVpzXvfi0tkWAcW5a23SfbUxKCe6MMXDtCM7kmm15kAa2fNRaVDNWYz+560NGjL3hs
gSGqEkTGMSbq7zOY5ADXLZDLeocNLSLKcU33tJ/gk7buQ0072Ekcnj7Lr391JICdvsLBYW4wlPBu
nZy3zyvkOZ0Bb+SeCIuGhSyWXX9r9ZJNMujRTtcwLaYioyOJxfPtoux3zy2gBl7jIj4KLVmC/BaZ
TyoPCDJS4CBUd3jcxPBB+ZieKBHrl2R8sK9kAhjEbbn1JL/Pcy9u9p5hffnJXjuZoMxT0QpMcxra
CXBUjiGsgSAu5cZ6DLwrbj8TvHKjNaD3gX9cyqAo1hsaY6yT/Ki4Ztx9kalBtnMkCold9jaWJ0rU
5+BGJuAfZvda0jEoTMvoRcwvNIBoR0W9M7bjE556N3A80DsFza35cEDGGSV+HZSX8VJY+2KlXRZI
O1wjqNyf50JYmPBCEICOz/GPBtwVMqCKC6a3HwSzQMT/5yjoiItTO+tHiAce0PqM7e66Itu1UxFL
8qqUcCSDBc0IfHnzW/xGPGbu6gnf3qXGtP4bEyVRoQq/hS/omKUaIBmA+fylWO8eHB/N+lVfAhwz
2fLT78eiB1IcdA1pLTmlLKffRAx5JG4UOZUGqNjMTBmnQWeiV/F6dpn8jrWE6ODTXh/XJuAL+fcD
Wuab2B8YcvZQUrPGuu6pxQjknSUzA1+iHBeS7eYWp0yAc+g0h6Xq9sFgsVrIF63vBXLtDTOz2DH2
h0zfd8teWZPXU1TsLtlK6Lk3PzgwViULeEo9aD15++R8FjsamX59/la27K2qdNjntoz1zjtXqUIh
PyjNymoNTF0iROAVhP71eAOVA1n/ofsbF6U9HFucjci1v2mYzL+Q9wpx4vYA8eA1DOueSSbBv7r6
iIvxxg8awv1n6pVWHA226djtGKsmrIf1DhTS32EdtyJaQAzSjLLY1pHs6/CW3FZAeTdfJ8X7qnwL
3mgILGzigeiy5MDha5FeXIaXrlBDQKzbA6EE29xiTyCkBPceDMAwXiMb7Qzrou8v+dSdGOW8oAiM
jr37RPGruwM5/wn6t9VVxWF3pToYcA2X0855Ddg6RBfz/6Db8I1Z3nacNhdjjKlpu1Z6R/0xDzgJ
AMSUowYr7BIT9glfZnOzuz1T9eMamaFI46JzGPmPrMbazKjv+vbJP6uNSiFeZu5Ra0W9OT3lHJLh
GhaolPHgT7DwC9CGR7t7t9QBe22P97apLWD6HGuZlrs5FJH+4M0r31vY/2wOm4rpxeoRMpXu2YNS
7gE9/b05V+mHVdaTpuPzy8qZzn25suhwq/07ZCpjiqJJrDOo+19Eb+L0t6Hmg9l6qQKtD/puzAwV
O0n+EiUs4cut02FX+wxOqCNEaBC2hRFjqWbMKRMjNGgiTyocGOd3AjZc1/bSB2OuvF80IgzEYL9s
TYDk3wdVazz4qYXpsOZZWpdYzXn9IiKtCDEOL3plWFhS3qa27oGCve+CLXYEif2bP0CjndTJbF+w
Rt4L6x2mxM5fb7cO3Y53yXLw5AADtt1MQ1ftSKvpf7BHkKQYnEidLRTja8b+MblizIPXp8bdBeOd
9UMzrZmqAHvwfsdj1xrwjNLhqI2otv+kU7m6JkI9lwbOtBhoawK8C5Kar7Q5CZ5NhEptftLpnnPt
iRikJSI4HlQy7WcRsTjB0RFwI4wJsq0xbXCTBoyEGA4JPI1wj7rHn//zCIp6IOUdIR8d3DREPMgT
A/bLI5f+osZW84VRX5hl4/0/kX+7lnVgsgc4dY9Xqc/LMjHtG34rGzgBFcP2iMgIBOeST2U9bkzu
ofUHNrozWErGdQLUvAUr5cOV1x3GkMKtati8XhyJTHiBXe4nuONESylvrdhdXBTpQXlu7xF8yyQr
IbJo0/5VgNvSbKwEvwBLumBM/dNn9gHgU/RvIa8uIVwHM9LOuNwKTQcB2/0+Ai4cJ0UknAVrUT/4
fLo/b8OOWNeOqBfbXxGLFyJ/MuFys56VTlNaiG4cWvH+Q66pCHNteTJ+Qaaa/3Zuear6EUBIstKn
VHK8QpfSHLm7F/lP0EZwpHoIQJ5O5iCzBxHkCw5GtaVRO1UGfRFblGEDKEr9CxlTYp+6QVyB3EQ0
TvLNvIQ8sGsODLy1JLuMUSYs9g/eRC56UamUiAXcEcNrwHkIDJBpAvCf38gLwPESeAwRnPzHFMDx
rAYxLBjHys3wNOpGJr1cwjsDHVnsGuAcuWopSce9h+9bqWjKbt/2/LmJii7HX0l2UujD2jXNynzC
0vKKGkV0T91YHV2Iz2ATR+M5SkrY7pUa96Dgg3g9mfGttPOTThctp9E6OulaLfnrGoxYDzmlYApz
/MIyPiqu6CKDt+YagIwaq1OsIiU8HItkio0T//JOOiWnWn0YCmWABeOqFNulymmYui5h8PLDatt2
0IZpobzTR8FZKNDtIQhECMc1QbtHBN2H1k5n+SuNMJNisMs/24eFvkucqX0h0j0R/xrxjxBZqifV
QFav5v9r1BxYibGnh7xDRsfXTjFMEQpvdlG6caKm4sIdUYGhVVIYEGwkJHj0oceT/bf2uQ7RAdcb
cB3Udfhgg9pNAG2K0Q/w3r7ukBTo8xBc5dpe439Q3J9qg3+wvoW6i0TbAnaxF8svKGhduxFzLpt8
4Lul3LZFQk6Uvas3L1AVAcfgbKnAVQWaq6idT4BjoHH+v6xevQe10ZDONwFVgmIq4D9ucqxOYQx4
DdtA2/fan5LOskGkYHJiZ1YSI18H0WMUHAzzRpXJQ9u+JVC/L7vqyyQptJbQVHMHqUqALTfaG2Js
QtyfKPqMN5GitVPxN6dGZt5TvDniszycEoD6DHSCVWTkSpJriav/Qbp/r3hxonicBLSMWmN8t7j0
E87fPnod+8+zAmJfxglJcpqm8vYfSK6EeSELvBLFoDhhTkiA7HQ/MlUrSSE9KPvmQqZ+ogiHy5OK
ATTTa8U9pebOHKBCOwf2ss5wqitMPkppXWf6QpEgTXPloGnWkvPyykjIY3st1W2DY1aazAndllQv
+a3fVf6t8n5LwB/OIRdc7xQQg/GSu5P15vqyBReVoSg0ZYCZYrvujZfILgGeYrX6HGb4W5NnZc4z
Q90oVUnnHM6S4laGwqDdjrwxp7NxbG4uJXev/+sXNR0B9zYWwt/uL9Y02oLywFTdkA5FkBv0TFvy
czvK98qWtJ+Us7ps22eoLYfKDrWgs4xj4ufr6LgYGMWQltXxXL9/ciC7gXVxvVVH8KjTgJR5LJ9U
AE5QI9/Gitzfzw6y1fa1hDBmZLZshgZL23jBvIWKLePJ8ousOih86ZAJrAJNRR4cOc1/AwASkifm
Ij/49Uhs7D5A7LGY19IutuYMNwxXe4ndAdcuGSGpDpRUXcfRoDv2zOFzg6MpF3qmlQpz6GWM5Y2C
C2/IOraOsTfDwx9ix2nHs7MYLEfLJeVBXGTnF7nAosce+VcLc6346UjdC8EjxoKfbbfRCciEzZZQ
E/MLVQIIpEvY/HzCE4J4wItusl7N4CA6vyyhU5tDxX6OTOxaWH7h59jLaXx21tUoszt63NUsIEMw
iVKxxHS8pH5bp46uy+QfybTZPR8oj7+OUCoeMfwZbHxT61ytFD92ZHY9Pz4FrbNIkTEh7PrpJxSd
493/1DbkZL7FbZKd5570gqDUpyVsdmwhwnbl2Hl5bEwpSX9G/He1/zPScpuFkZ0Xyj01IBrkAUz5
vB3+KYVU7D2jEP+zjIEv2KC8tDpWJ70d2E5VditIT7/AAcjOWbSonnxB6v3DXnVwoybB5RXXHH1N
nN6vQsuEF6rtAiF1zivfyP69zJSndzrtZz5tHbioUgPkA8MjiryAgtVDJI6HhqUSvDnoVVuCJV1F
WRLpZI7r5PJcYVjMsYbtjaXPhWy/NWA2oXWpqNAiFr69OhPaZKaHFBRcJJRBzzr1MOQiLTGHgtIR
eblzqOYAj693R5fRgvj3BtKOtDKxMILFfGJYjsD4Om86LcnYFrrWys7rHNP7Ob/qif4kzHusjVnM
PIF/ANZUVMGCPDt2A0pIZdoAP8Gc27oDpUFxk/oZNVIldiAob5VESWtuxFrTrZrtRyqWkx4/MrC9
0tERIIy7QojGFDIOmWoi20F/jkwpLFPncq8ODX8gIYMTGoUgle7VWEFxI6x54EArQ8w9MVU5NLeL
PzCFQyTl056Q8dkuro7Vp5RKJN1y+tMU1N+ttoRJMPSb8GNjGhWZeCsfgMPWYjvf7ajs5Y7xCi1b
spDRKit7IBIFcaWShYL1fxGfyF/s8ssZbYeNcjgall9FqY5/qCAE8fGn/1L/oSTwU76R6DmfBTTR
tHvXlTkpyi+68fDZvYGas6fOUufR9xrlEAysQ8cmTmIyo82sOaIVkxXrrHXny3JMHvk1uvFTQpAo
+2bQpVaLoFBoulg7VCiP1woL5gyiq8sFHEwWLJKYp90RKvaI7aF/T85tyI7agU2hJdElfyQ0u0dO
dg4rk+JQ5OWorjlsL188Os0ag4QE3kTEoNHPTOPuyf8frZIKGFoC8xINGVh5IID0F3v/tJxauUyh
K9RUyAR2eUa/BIB1nNiqj/S9iG58oCm3D4wR+5KCZeAuKH1cMAlRKykuSaLgrvojfOJ3FD7Z/SdV
cPRv6Lje5vwZG5PQdDKobhJOJMjn9Dvj6TqtF1jdMQOTrBMA7TVtz5ZWrMsl7lbGI6l8LfKV9W7d
wcDd8x8+ZDCUP9RB5PJ/6qiHzQFhaVFLptz0jqqLpfmmE6tyX5YuUnnqfB4xmvP0PGf5+DMYwrfC
5ZPEDKqBRrYTkp3CBj8b3iI8yjlBiwEYu70DI9JeuWuVk4nxz+QFD+cC1VM5zid3u+PV6wuXOZuL
/u2O57gaHVd2GPo5nzzL4sbclhG7cX2wNing2g2sXf4HZs3apc/PLSkcdamXQ3R7reNjGwMHi1ha
jH3v5fSoTDu+3tXnTll9bQXHeLp3px0DNujlN6IUL/2CsP1ZEsl+6Cy9OyXSTvpFuxYxtRLeFjxs
uLiuftB2Oc1rdBfYxexzDGIVwbJ1WXL3rngdn/gjm8kWffPmzpoGhrnNh6xBhLEAi49vvjSFuIrk
lUtSH6M/D4iraEQq3d2kViHNNnpXDRdcaxukxNl4Zg4HV0D7qdsleMmzUdYu1Gv2gb4CYcCPjDFd
FqKgOGbtkrSkU9BVhU59bnEGiImXJr1zTwoEzDUWuxc9FDnRFJDc92doakVUptKoRP+fzAYqYYK0
LSymY3Kxyn/5nE+jNgT3Gx3kk1irBJKXapPMsrgip/iNmKu7QBPAXDggGjrGbnixkUkpSkCksFJM
boSFN/CfZaSZrQS3yCiPi8xAMQuJbzihgoIM9LGop2OSGGQg2qAXwMr60H8mldHVqBzyO+K72ER1
0ZzWCnZbClHOh7ZCBQWHxzKKUkroLDZEnYZwya6xi21o6re/wR1jGL6MmQpEsuAH84EKs6Q56M+U
rNw77Fx52BV1qXjXrrH95EEatcgkVw5+j6EqdVJLgKPfXkYNvGQdfZ57cpygwBu4dLxXMX1o++vi
WM5G5z4YUbobyl5ajNGebrDNQTBQfD99JokcRwzqXTZCk/gZaMscQChYgmUbNrGXb7SnKL3OI+me
tLzUfP18ZU54hkOX0ux14jlbftOz9FbHCBW++WneOstAmzsR/mXTeEfzZ24i2yUu9AGDlvicjjw0
JanDZLaIhkXQTnrzsdX5QQrMeO5PCTVZeoBZNUiJhqWEFjnv23Q/+2/tazvyjbS9LqxkP5oSiY4I
aMlvYmw8it7HXfdL6+LtAOiWbOc5VATVcLmJbN//GgQ6NIz+In7DJPbXppz9305bxiIzeH4kiu/a
Q2AirclicRZevIooKgAwu8fvKgYSQQOLVWg1OTSA4/dlfpWJaV4mjXsV40pZe8yDpGhhdPNwBT4W
0v8U66CJ0SqHvmCMKz4PUP+SFinrt7ENN5/xRlCjSshPkCYeg7slZKtyw+nmdKg899Y+F8uou6CH
Q3eEkxUhQqyDs7Es6HX3fMmJ3rS6ND+CvNXt1V3/qWcbhAsQQ7o6NakrKsHojApnuqX93o2bvuX3
A3eQF/5xB5xYm4hpRUnofmuEj0YtH2EKtisZcb2rDbwq4BzWFkjmiiQPruun6fh3LcnnxDh+9Uas
X2KRAiLWWw6Tl2iUPTpR4sJwylGDsyJSEIMwD4w+AFkscnrh5a7J0rg2LaorUxA9nNeewSuOdbOM
YGQiQfbYBCfIW42Tz9KvVf/heJANd2xpRF2rp9vb0313dywm59I0vajF6X9UotK6/KsawmTzlPSH
Sj0zQXts4YzmbYkMRGcoaZTW7AlKwE2OAb9srHUZqpupCMr7nfqQukduOW/qOqjz/okN0aiQcT5X
MR5tiIcb9EGBJK2jyl3Nowyz8H4hmK+ZobaKiCO/PXzmvzyvehJtyahBUwqGo2AdT9cg/l2YS72f
NJE7Z2pgwHflbLvQIEl/rqeyG4yySoXj+Wgyz4qZbzyHC4zyZIBjqi14imhLFDGc+3zMWaA4sMlj
eFrr0JaAPqR3tQYlFsCnaDU03mbxip4Ch6V+HiiaNgOEHz1bOTMQOPzn/pDTQRCVsHCEWIGwstB0
wl4HbgvgPBuvMvRpug90RJLx6dV9fZs0VPZjN60BuX6dmmR1ecYrs5JC4aiC6vi0BblebEVdJx5t
A8N6QzV202EA8tueLhHiCfjqilzlStGdc37PX9xMxe70qhYhvnLN9F/graAc66tA1R76DydRNXHG
FHVklsrl2qINTKeynpPLOJfvKyCokuLf3ilsk8L0+IeU7QBfwg/rTZV6P3FXNsWlS+eayGRzREJf
hpCTM7uQ05LpfMdv3/mwvLclj108SLpKh/bW7KrvP7ERaEkKzFgburn0NPbE2C2U5gIoJtDW+i9S
ooisd5+ceXomqzkQVAdtAIg+N+xzn+0+xU2uLGBlyEjDuVbgpBSk/qQwMD4gGyWagqz7Lv7UUcum
KLqPKSID0meHoOUX2MTh7lFFsTBryJ88A91Q8YVYywvbJnh6bbfpzbNZILjkYoD/chC4+v44/Bct
fstzAq7Vg7V0D8GkqAcK/44+mOHR+0K4WOnRro2ygJZpb48n5Z1s6Zml15XdmlNPA56GbbGJROo5
sAn4/h3jO/BGelWV3p6C5Lt2GMkLkSqioSuisf3c6QQ/nr0+x9T5/aQvyXqCnORmpWE0FrKPxKmL
1kJOuhr6R/7VpQWGihuUEWXR+ZKJkHd6WnyNyQvInbcBqtgNOMfZkiu+fzGyBsTBHBW2IwjK9E93
A2LCyuEtvArlQVi7/Fs5nV8IFu1bbfr/6/UamAEV0vrcNI5clYYbplnjc61gtZqrM7HbJ27jWc2T
ysBvvxCyF3H+JPTbzm8bfsq3j8/Axv2+bMfGn7RkvkwAffM/s/F32AF/B274YPLUUeREw8cUQaJV
SALgF5ybwMaxyvnNCLoLPrJDNyXb/dZD0XHTtf/1762OarQBW3Rhg1UUIK98uVWdjvJzDqUKfcQn
EYKLzZYV+x2kys/OqJtQT00UCYmNDSNZANA0+3RbYK55ROki0h880KXLCPuoX7WIcoV/6BCkMigq
Mi3xQQGCtFl9gHmRsA/mGWFLB6ktjsjgxPCeOCmYdrz6gRnZ8DrHT9BB6wMPj4tbqAkvYNXgBJjq
I99g/bQNhSlz/KbpV599SmPxXeaVa1qYbj9mSHaBtaTIE08dipbTQu453hSgZ403F4h0gnJlLILs
mX+Gak970wz0WDmGCnOA9DGSqkEzZPzebTDSOufieRjIk8wv7vAxxW3BSGdJhMWZ8ZAtCnLgh2om
ZwjND6Ir6CAYGixjAZbNeiSJamF3AQvV5uNQW6BrgXakW6eWnQS0DPb3NdCvFYYVd+f6d77+elJe
ybrPFxVfpWJdumsTOQaa+pHgeS2rmbToe48XxT5K3noVAvlXkFbGcOUVeOW3aBNksTssd7zRmK1g
dPmG7lMcB4vqzNw7ubXhW/uZEzLdty2IZqLkOiDKndqbF4EUjXflvMxtM4LlBRwbY4MC8FgzYoAy
yL9d0ZCtc+IzCT/jsFbCcKF7Er+mCD79HZp5eeW0jbYz0SZkNMMt8FVFLVNtVqDP23AeAZxeXiSD
06/l06fsjFgsG65OXAh1wpelXrBkgHCgVCnV/7L77hnw4FCeD5Y+zWefA5V/r85ZCRr5AQpt2nCm
9IF04zMjwydjNinE4bIeV8n1gp3+TbWNGvWm1twOdJJXrlevTN8mmsKywbJq7AAR99msHjdL3dJ8
yrnJuRaQGjvvpkBdt51yDt+un/bZV+jKtwMpQUytDDUfmkZLsT5mSfEH+bY7OL6lV5NuDrJB+fDq
XJAC61HbbSaHgKAv9oUmJo9DTng7zdYNYjeaTOEs1bY4uMJFki9dkbcF0ElxR7o+z0mBquB8iRd3
ZWc27GVbpODiwQ2iZtEgUzMUryXEXLD/DGKIk5KH0qf2D1d1wgbQFnD/siGy9OTKGy4Efi1DAKKo
Bn16l+z3U+yS/Wt/GC1sPhvS90tvoZcCEGprOSY1HM3Uge4b0l3JtCACNb46fwU/a0zvl5eO5fq5
qEFeZW9bc+bmIbecU42eHgDWKkA+HOOEohCadTc+o9PfDzhUe1IUys2fZvIh7pQPO9znO85IS//9
h3K8VWGU3WL4nCu0BES5qxJbjEOqkANeKhjhB8SCPjcB3D/B5R5BoSdALOnzadgO8/PCMRnIvdEd
NLKO6XlCVZDTgGxpG4aPgNoUkWv/tzODJkqHl6V1sj//yendBqjCADjL6u5rMOc5MDv3fqAG43YQ
Bm8sCupKWeqdvUVlh/uhYx4yoxpvhgvSIm4rNlqedBYTnuYZwqk/WnocuCNeOhEyOrdGy4sCLoBa
NLNQGyPisawiYkeR5aFUjumLjL/A2e4HYR5t8AQviWcPzdSb/xYDiQf0pl47oyxrUV+Zx98SM+qf
QIc2D7OIIolWYYu06XKEITEw2JRaCsoGZdB0Au53ffX3BLlamojRvxW/n92nZGYNIYB4RPfu/vjM
pI52PHzkKa+MMjddXmeEbs9pXAUiBbB47oGf9Es2qPCw/+YhIiIbdhoT352X8Kn9r5/pFFDV/3G+
o8JyuNlCDap4FuA2JiLoaLrvkoExodFXbfrsK7Iq2KrWQE+AJsaWftz14cWUolNsI7TMCDqd0V2S
G1DJzfO9c0klptjbMJMscjHqGodx8a7mbyg5cE5tqrmLN/Hl++bdu1jXWOkqie+GqG1N7U1Ko+jm
JYOsZ4G6Jh22QW6roekuX3xsXNyWC94i9l6iR/7cOAVDaALrcrIRhDnaE1BHhmcpma1dWb8r6xLU
9apBy2JRsZhEUnHMVwPXdxMgzkjxfrGzRlPudud9uiEsA81zByTL2kD+26PMThldAl6371emSCxa
Q+7yqQcPIXicS6a2wXo4Wjc2HcYX7yMH14250Dx9J5ACgWfMgptVojHabjyxYvwvMT7sGQ9xMu9p
boIea9vAkMOyztDrJ17GsNeg+dnJAU/fimWPeIHUhY4R9w18Ck5gkFEFgApZOhjoPhnZsy1VhW0/
GMeke7B/NqwrzyOWM7BNAOSX2jDb6Hu/7ioA7KXImIeB7n0mYQuWxUnTmhEDYsennjGADdHNpZG0
JBrPYM9XLYvYaiPpv2TT6+F9VxrvFFQzSfbkKkEMBWHwqwE7KOB5dLCl4Ucpiq8IEEdCwqxlXY4D
rcTD7bqkU4270I1x3xrM/ASSE7WpSN5ISzMcl2pEkFNFPud3Sj/hDThqbh38I5rgG9YOLUCwesSv
UndZdv8dZfb477Jbm2TPaszeva4fd2zkQmcUaTbgXVPcIeVk0FOlNP5yiohWcR0Uh4TPpwvVOgIZ
vpZBwil01QIe8CHULePHW18SwhA86IapIvOOE7zoc98FikLE1Tkj9AjG0s/KmU3uB2kuQE67IKkd
tkqrmeo3BbZ8V7APalx4G8MFBhMathRHnSLX+oZrNLXz4cjdvlR0jqDwchu08JiHXezJVucuZITm
ubeyHqL8V5YUuFH++j1lC9aMDs+M7PJw74uQHAybdquTTX3vQ5a9Oejz2P6isGSAwsNT+Fn3ds1T
xKNOheGdVo1wY/wF0BhJMRMw8DBAo910R9QidwEE6/XSL4ZQRSGqBI5w0xvwJ95tp5g6oSva6JPY
x15D+HeBfGIHRt/2QW1/W2WtS4PiJopTaID/TPCovNaRohiDbAmMwaivszXdQIvBr/OweqkML44i
wUT7SbbfE7i7aNfmdJsu35McNlJqrOch9knTTXSlqEpflyZqgvqRrAyCmzbFYeKDIgmy/BjOO4kW
PpdX+ODLt2uf4w4EeZnFr/8QZdO7zU02e4P0jKz4yw7KY6Iy/JX0SWhZ66SOD4BxGdbHkpNYGM1J
UJGBW1nJj88sZ9bToPP19mEbCu0WHcvOVT0pUk5kDuI6X3w0Ma2aSLfXozVRUd/NdwzVqSi61N8q
vuohJL/8vGkY6yuTag6Sn9Nh1IVRMW+gUgDqNwskrSt+zeUhbtNhDHVEWXKxdW6XJwUADnfmcwJs
/gAbUOFhuZssW6EKm60ywLoXFaQMrnvHVXiirRaOrwv4IT8i4ebTslKrMNpXYM48XzvCfgA2I06o
ZU8Sx6uADp9NxurBBRir03YMDrscnF5hAETNebxLe1I9LNsX1Tmg8i+f95owLd/Jh2nLCJW76cpJ
mbCg5l8wdZiqGLKFs9A3/m+WuNxx7qrjOZ7dXBaLGcNnoe/GXKQ7gvkTda+p0i998JjO8i7zUuJV
qNr9s5ljBajKt7UFrs7vT2Yekhn1LS3BZUhGBPPekcHbqYiuf1f/mGU7KawSCWJG78tDkawvMoHr
YyCXsigNP7gpld+e66485Pn1fkEBtXXSxWjNpS+FpL71mVk2lKYlOHFx/9IstyA3Az5cEhFsyxzv
eEBsYsPP/Efh0n/uUSL39CkoRGVYoyRUErIrLQUEzxJY9js2u5YCJoja5YjSwb6wiFd1ef3afbtf
2KplJ0mNbKnkasYIfMCyHVY7zRd5MQenwKT1pFlEkC6eKT6DE1VFpcpdZNbbC1ZyVdJpWb1lczPi
v3Ge7ixcuN1oqs2007ASJlX6vLa68P0PG83d7mtfEaQigsuOkQTGTePAj2r++CLswV7bJ7Wlqvvm
hfdqvXqrnU+3FxYBm66ybJRX3wtOysCFhgSdmQ37y/PoCVz8LlOMSYyfVCyyS7pT91Vh8h/ZV+jg
35MlJ1FaJxatODS+glxMKuki9VElQ7vxvVqlHNq+1A4LFQfBwqxDOHRK9jHihxu6/W2OVeL266e0
RsZ385NTZ+F7P9vUkY7+GQ/sEvoOn2czr8rZHb2YDTPix+7Uwpz2hQDoHHRE+2zdRqHb7odtl+x7
bq8v4KUF3FaXDHYT44VCbYXYTKHjX+H6uy/5hWzTZhUcYMi7Nhhns22EcXkybyb/5IzDP4QXC5Kc
/Czvkdtuqjq+iRabnbNuv3DQT7gEHJIS7l8Myd8XUFan0uqvBJSf6DyR2wsZ24YX06Z/L4FS5r5o
Gvp3KlE+48k9NYWeQxmjtG0Hec2AJSTIVZTQkcti3xg61NQ3hnMmPzIWCEeNmwThc1VjD0VpyeL2
3nzlVt2/z0htvlq/UgApB5qqJDN8k1E9D9cCdiCyJOYZ+pJxYEmo90ZSnkckXJrzOcGs+od/d0cW
dGGGFfJmtpVoly6gesQYOnHU4FFRc4OHZHO1BBLDYtwSuCfpV94Ma9KRb8bzpUFAX5XDz1TPCZs/
ANUT7KxQ6zsfTCfkk/yq5Cb8wJM3RJ4dxPB+XCwEm2/ivmYAlfW4DKDgjWJtAONynd2Fu7lwVniu
AicVl0DZRsV/DAWOgMtufFKkjFxnbzqxpsk/UP6Y9ayyP060SmpGyywZYojWoNUGO/2Q4keh66Bz
6FKKicQ/gK6F070AbFsz1c0cNpwAPVJn1nNruqOeOvKe8bgPOQWUEk8CWIvzCW4AC1VPu2q7nsyZ
aeZuv42h1FFqu6Inkxol+8UJZE9TtS38DHGm7WsnhitQfU9hOOGKl6Lz2uR660zKPCp5zZyb2/JP
GSGld52XCmD19vmCiOhdnDt0+PUix+cFy1sljo1KR1WUBkmIfCCvKY3fi25Ys1XxOR55Vo1sUphs
sj7w1Vs9nnvrNZmRMbymdpbm8sNyURO3ayoE+gxzOgO2AqrcN+7euOfcAKFK5keMGoksh/DNM5pS
YbLuNY/aJwlGP8tG+mg4nMzicRlXPy5jMOc9LahZiOZbm2pgbtxAEhSl+namYwhLeYww9XvzzgDe
9Mgu3VebG28CB8M6ln7tBqZG48b0TP3GEwATMY35KsoRye3AunDUZcVyayu4iVmRhibISsRfI+SO
Is60IBGP/GbRX80MkixPLDhIdbMG7tnLd6cS4X2nw9RtNJZ63OjQ1zlzjEH3B9ISpKWyu29dxeDg
6wSIDFZpxnAUCpwBFIOzjP1dEsS91hElsRYTvv2VU4T1QjmrOqc0vwm/Ma+/tgVgVVYVDPxTrV7v
Y6fxx+fv5a/BuISLMCPkwyrqEYE7qoiDWsQgOfryI2tQrOyLVxb5NagkFB0oA80tMFnwXE5ttHKV
14/FKA0id6/Z53AgqI2h2TFin0laVmV9XuBdNGbw/PzVRfrHLPewNEMHkfl8ns4ehXcNQj84NyU9
KAn8gaKjuYV5SksJOAN/3Zm88F8uKhHbSMDyoyu5ZTOvixIqukYI+6pM1gwfKsTbbLpe3RcPwzE0
LJ7UmfiKGPwJR7RmosK1XBS5T5UXLttixgD0+5fk3shVnj3c+qnFoj3N7dI2hf4R7oNPZZjJUJu9
R4pqPP0VK0131g4gwDqtzgeaUe5dH5Q451ZmFMMGOkCnxW8oVpydpEsdBkIOVedx0G9aWWCCCt04
2WiThiNhbr2bKQ/XoN2R2PgC1f4iV28u8zz3rtPrbAiocTxgNH8glGyPX41obsmkshYJ3+73Vcb1
Lz9lUS2kb2yyv8Ntsw0aV8b/m6MlXXcBaNCl6jRPtk34UVlfb3Hv22CHTmMrZlUiLb6t0u4RbkLk
mpmExL8MtoNsjFLs8xQtkZAt9lKszK6qnEiFndfgp9YCJVhRU0fdwk61TrEr6SIJjE3NKTdnjz2U
HwnoF2X8Y7AmFEdXoS0kTYUzXvl6gTmGisqZOLUnP6sKo1jU4LaxCW7cxnhmJkSa16UND6aVB/LS
WFUy+grZZO8tlieXOzL6quH0/5veu14BleYf8OhlNOpKCWyZ37ey56+zVnOldDAnRIyzvRaL5UKj
T+seX415d5irUyFgMG3PYisqvzMAb/Wkpn3gjpikfxxIxmtCmZNtguBrLi+4I+SAKOaq+Y0nnkLH
lLETdn+H8CnE4jMHazoimyXDg0kyw6n/uQhnxWPvUaVhZbGjh2ojp8zZonPfCm74FImEx0W4tCZd
OCL04VR39F2aRD5vkSCB9pNLrKK0soN+GkRcA7lq5qVQEfy2ISJh2FYGit/mEa+wxPqywl6nRPpu
yLUG/tfVNACRVcHrAMXtR4TLTYmP1bmf1HBiukqgkc9LJR0zG5UQd0pDWQfyfK/utuZo3L65J4EP
pzKMWSS/OtSU31UxTONBy8t71ExMbTRyeOz9lK1iBufxivW/9eFj7RcQlRyTZgY3Nw4mbqmQ34PE
sbMbsSK1IYE/iM/N9+YXFi6QHyuUnrjBQhR6halXKApZMdEZboERO5hup79Jn0O64sQJKa+Ut078
Xr0uAk7d26uA5J4pCpVQYqAMmCPqIIUrAhCuSgwaKGQv8gvm7uAMgsOS2LN9CzuDzC/Mop8Zyj7M
D01CWhT4iAxyNanlgBBfbMPA/+6BqoyUEYj0ed62KsKy8WTecHGKXLVh3XUHIjWfu4+o2WNVISTR
aXoRGKrXtuY/bO029KeQYAcnDMbZ04nibWEKPePoF7Z4EmAeK/AzUCf2LGrwqrAmZCoZBNrARqOp
QBrbOR3O3tu6X0OFVlUHCkHOQ3W/ir7UZgyZhgTQ7GjQCXTXzcPX5/Honp2GKwcmxrYzI7HX86ef
pZi8OORtLGkqW4QuZpObgQ7KuAniDwlo94HJs0DT39BF/V7c4OAj26JiBW9RbImxvG8ufOu5AW8S
OYKumubMehjeWxLODubZ9TkfavwDJosAk935f06iLYxxqOJow2lcqe4RV3IshLD8G2b/ORwscad2
fgvpSLv/oY2X2xXDib687C7FtTajtEd84HrxKvReC/w/GEHqQiA5kIcL85je1UBLvidxzEkXCOgJ
cSwanh0vE0/vtRfpMMwuqZtjM6dMFrQGpSmHYCVXlA3h0rRfoutsMLF8M93gGgXBU4ZqFGnbI/FB
mwojFuy2nrwiOqFJt3Z4z0ALyjPa7zMt4PVcO8ldkxmdVceWCjR5cw6PYDhI93snwjB62lMCnZOz
Z3YvFPRgfCkFMh91o2lkVl8G94FQ+W3PVhKR7K5KzHYQ9hanzoNfDgiNoDULGE8sBEw46vMTVs1V
Hu59Z+Q40+vrVQUHWpZERL63JIrHpeO6qBHR1wxDr0juBIURaUIw1UKZT3FIV2b1HCzOl8YKc4Lt
/2WCedqMdOkRV6qh1e2swx4F0KewF5p3H1C/TIMCoxkFhDuJGWdudRdMf04UObNp4flZokYNLkho
dcLC+nBZ6eEshgpG7B4BW8yipAB/K5Es734cxpx3njqebKxDY+gn/a+SbwQUvCMnpt9IjtJgUiuo
+3KqADnxTOkBytSc8mjtObnHkjGoBavJ4CGtLT5Rn+89hxCc/VrOWe+x2S912jbrdtgPkxUKgyq+
c4N8+t4fkMSdz+LFxKo01k+MD16Pm8URFZBHrBXr/w/uwvU3NOuE4VDUX+QQqoFz9kP72gZqnmHC
lmZYDKffIBLX9gi2UVnaS4IBxxzDgoc1BvriLSL+7VdGdLy9qTfnhUrkCpON2T8jFP3B5uEhXrC5
BnA3jOyfClnSucW1uwj3tf2LRBWJYce6BI7JQia4PotGegmebQd6fxU4roj9Zh6Qdd9OnNnfqqY5
WH6TRFI/DowBBI7fSk1g74Fyu6soN7AAou2zXdOlKTUylvZtYMfxD0JkLGrxQrZTQFalS2gX+GQx
Rt3YaX6v99ND08ErdCvf7yzs02LHxx9rzHCYfwEATa94KL2Ea+x60IE1TwO38Nzvl1xB9ALLhf6A
IWtu2GhzE9Oijrh6wUvqQ1coM9fBqTamGPzziArTTli3tbL3BXsDvDPDOz2PBVdI9dHURljDYBL0
FOUKtrTvwf7teBCXmGpJYGc6CZL7tkw5+U+vwX3Ak0oaVeVtromXqsmDJAKvXLB6ew+zX737cetm
CCDhjpF5vw3UR4+U+AQmhR8Te0V48ITrXHrK0BN/QgGjayzyVOjfeN/uuyU5f3E6fo4xxB4TF/6u
jrxnSxgqn/vmsiZN3wh5DnpgCw/WLFgX87dqBoCrzuEUZAvl7UtRePZeDRrITMI/vy9YoE+ifJOv
A3yhq7lNiP+i8Ye6OTmVnTugVDfJkGVr3k3bys5CKU34/MuThPLMzRoxeUO1EBKsTo92vKRlfmFk
wykncZ0LbZq/Ali2Wrb/Z1EX19yMrB7BMNJxYO3fSn9SYdQFnj5vrs44pOnxzcju+ZdR+YjuLuC1
buG6SRCjABCImYONrZ793qlLW6IjA5BW2gAPLznSuv2Jbu5UGVA15EkpqDnB8UM/N+BzOnQ0/Vzy
hq/l3aiJZu/CDpLdkBlDtiqQKnNHJqnQ5id0QrCbWv5Q1pkx/qqwCLWLNLdTBJ70FkI4VmkxURYh
MtIOUJEREbzLy7v7o/MVG2aKxrE6JjJLTjphKr2HXw0zao/ZIJo+MrdEUqYshDgRIbIHK+LJVHj3
dHau7TiSb1czwq6EFizOFB6pfZkT77EV2eRe5npYIU9Gs7tWz0Nz08lLJ28TNu8GHaAQHxEMktpa
sX3qAMtActfrCE9PNM2CGwrCHh6lTLowop0Tuy1qqQYAivyDTKeqQI1+7okBa8JS2foKIN3ctwjX
OBUrc54ldM53oG6Lr5tCrvIz1AtiGnC+QGo7UmkpBDE0rbjwJqF+SaI5TiJlMN7Dsq40bWxnakTr
1Acyk39NCgow0snrwh3u4CQyQU8MsNF4k4OMLzEHuVoOXXrhikFi/cvFOKrYhNUh3P0qPb8xR7td
OXeZSTU00ekofOYl2oR7G03Npq6q2J2vYkdm3O0AibCVTQXY22ZJiBkOK8x+fZx5DmhX6IDpClIb
ykLkVk2X2We3WxUn1osdkIMaXyPLs1uqtkea6t0v1yZn4nN1vq9O/B7byJzTiLodDyXuM/g2sAdK
wz6Bp+1goBqkmDSsmEdR8C1pB2d1PBt+Jg4dwpmr7qadZjTOZt4/a/dFrl/GvVATS4pzRjakT9rk
smr6LeBWPwHnilUDwTo6U95NcQrkIfs/cP6fgS1wchu5GHifJQ+KxUbR8P0igsAKVOIRjZP+hcVz
wkcwDSdNKpaXAPZYBkyEdnZ3ZwrW3jqsbw0WtOPhRSURXd5IlEwos1iOSpwWuybUeSHpvTIcT3Q9
sC6Xvf0Vr+QxAbKcUdjiWR3JK+5UP9yaP6522YoDqWMwUmQwNsBplZLFuhOLei/amHH6YjxhjYu8
c77M4nhDNUpS23RskFfRwGfsDBP5pbs/mqy3fooPPIfFVzPUL+rP0jUvGwxDy7I+aOCMnAL9WIQc
zN6BpJC2tzPenAoOVn+es58qns6oF2b6txh1wsUyTTEwO7FXAXfIEILfjdw9TDtb34P9Bvf6PxxJ
95ZQDL+pY2inPMN4g3yjiePScz/Sa6Q/fkPJLaM9CAAYTPrxMJxryTCTzku3ak2Tiw+1gVK4ZnjK
8WnL7SWFUCiNftgE5PsHdkmmDqer8AqjMu3Hy2t+Cbo36I5bsNIMiJKmjOY2uUwcRTG4wX0cTJbR
SaX++8nSfcrJcqZXuGroV/47ys8P1ndgXJPKGV/R+QNsjWaujxr4Wc+zexAsQEWnn+yO1YjsL8TR
6tXYZB91XRC39Wtco9uOWWuWKtJKVoeuSNQ+2CqT90iKWd9OEApfEmVYx63OjIvCpawgzCt2NiIN
fEOONqayA3WMRhsJ+uxSL+0Vm0BHWBftUHVhQrxU8igHlqzACPkNr3FT8hd2UoAsr6RzuykKAryb
tyJeXtBJ6oT1Rnp3QSNGTpr5YkWZIXnyeblKZJjB1N8KnFlQAHHFQ3yJroqifr+vvFSon/+xbXkL
6gUb9/w3vvPt+IwF0H/6RD3CPrehOEjixE6r/MU67zT63WkzrgZzyy2N/9UXnouItOjShXimIE2q
OW3iRvMKfpjQ1y3qAjwac0QDxvtUNiClnNjpZIhtSWFvk9+KUVTbxQjW+f0+RgPXQoVSGtq9eH2U
dnN2/devlnoAgwt/fPdAhTdgjrKXzAnjszfrAVyYcHY0yV4Qb1xAjhJy/yqDYhQL5JsLxyiQcLH6
6fFd4YwjpZ4oFyMQICmW81puhin4FKaCHKc+pRWdt4ee4kob0vLoZ5KUz1cXuZlzgkYoRfnfFKkR
M0NCfL6JuqVKjB1zIZCBgxFmUXP0Gu86GRHehq8/BN24pzuXd8B8IRKg07DUaw0NaoC59TLOH4/u
EfD5I8+IkvC3RFOZC4PC5GVMYmS7M1c06MAd4w06LFc4ugOnTwxTmtA3AOHMaOrMHsv6kME3FHeB
fMFLpj5pXTpy28jIenTv/E8XrGoikctG1if9yfSY+mGNB/8aCfwl1W8iIbjvthLCoKgll2lgtzcT
r7ZljkJ/xbPiGSxc39vYtBgZ44PaKai/hur6kBDxnkaQu7x0+kIIlouye3egtzKsKA8O+dxUwOHv
6b1PPIb32SxV2A42AAdys6NijeWUU/AqjPhOUei0jjI4xiWnIX2uhOZRJPUwvXNX7lBW1HVBpMhW
16DDzRI8OtyOBTuEmgJ+jtIciv6zkcGAkwVeDdh6A5iSQBmf20JDDgwmEtbfIebNQwiiajdiqoa6
CX/uCAyEPuWQF42vNbrAu/B0tXR97nVfq7h1pf+jyciI5sJVWnEBsL95hqT8hIrKTDtavZhse4pm
viNS/Hcl2UtDBnU6BJ43gLXy8Qqy3+VvZX0DT7NaCf1jk2fXwsCq6Tpy19nEKBn3p/EE8dwJu1IA
QPKz2k1mSDxaGhQspFU4eDsNqBKo5VZ1kNuJGODiOQi6uLksU2nr2CEN8s+KRtHApivGMEd0KPTr
0FdAvWO+lPY3sno+IUhL3Ev/R0Rua1fmA9ritgC/8toVr2riysJ/NfgKbp5uKsnSY9sfpZc2tVas
c0ceSSXXBm/Dw99gHnE3lj7ZEutn6wqL0CVZc9p5IB77Hx9cQIsc/kGiDfMoxm+yY/CxXbif2/pk
l71btcaRnaLhGOQ7RnKrOuAE3u+tjzoshSB2gW42UfPBFQRIk8x4+RW10bHt417mz1nuDMEl1Cwx
BCFO35bjNSA88ZAHvF4qG9Z6eSsfAQSuzhpNTa7yuPhHeMss3AJQGz7CYv1dbO273wG4eav4SuK6
9GyTTPFY14Iztr+1CMpaTcUCSAMN2gUadOp2BppSCB/1CO5Ty/BH+D3P5BvwDq3tR9L3+9l63nrU
FynQiD1sTcGB64rqxZfCH/Yca5RX4Bq6i4UK+N63ao06p+dy04NXzbbtkDBRinaPQck0zijcscBY
9hRXPMVQo+QWi2mh2UDIpXcKwcR0i79/K7HqTYMTT4DJEpRyIGyieqiy5ZPxb0wefadRVgM4O+lm
XsqHATtocG7Qz7OxqaP8FbaH9MV+qAPjIOhZkOUfyEG+crahOD5Q3v4Ab4MqgGrML00yXSlG9IwL
5KLJCXeJ2r43waFHyErCE1pyI40ORzI7BcFVZfN7gYd04RPcc3j3BdinfGXnohq3eqdiiLbheEOL
0B7onrOUUjMxVllK1BI88dj7xGqaOgAcFwkqex6y/Oj9PXIaGKRVH3A5b9ssdhnkSo3wXfmPqj6z
rqat8VKkwtdLIoJ65IuNe+s3H0vsmoPEwr9lh/DQCDEzCwJ25Qh5Nsajx9c6ei3sO8SfK3M2CLCY
aEMCXi4QCAezWCPb6r9dh44O3VuW0YD5QLDPzaK0UOQtLh267dgyOPf9UIQqIxil3/VwpQTcgWEK
sSxUvporEXLeMG5gSDgkihFlNfV7JdL0F1ObDeKJR5sIYlqaPlHknnk1tqrfCfuw6ujtnOmQsfum
7QbWXdrDWPF34SBF12Gb/MxJ58byAp17NSWhy/qB6Vzzf+ykLqqwE8waY11iu8xQW/jElNO/EeHz
zaFC9o9gTMVYHkNYujzPrWTygZqqZBxNM1killdWNFHRph2saNCq8CtIkOzL7gKUk9xYtcu9Hnhp
NU6KJeo0JvctzZKtpoRpvV59BzQgS3xphU16a4dafqJmLmhpv8DnozLBBsCJ6ol9gKDJNSUf8Fy7
I8Y4KCGH0f4mPkoswYfLZf7NpJEpGCxqKW6AlPQtZcLh4+kWCU4rK4apMag99hBATTrWTpbft1sQ
W3qT2J10l6WUh/CnEpcCHjpluIdPNQSv0bgic0o0Ev+7p3NoKHwmvtw7F1KQtGbp6YttToVXjA0M
1wmXhdVNGLS9opYHGCg99uCYZm7zgeD1lLCgBI46EF3dLqzIhRqj5MdBUvY00i9ZC0nk6z+7UVHq
CmQ+rzAJkr7OAxE/02pGGIS5J7X+6vz9h8by96m/VRXjRcC9fg/mqaHAvePMAFUUkClXFONw+j9V
YCa+rZOtk0nA7zQ6u7Yg8x+HyCOM6kHh/8FgP4nM4oYpqtLJYHNlcWLFMcSdDgWGD21xv/S09Kd4
cooFa7XaHE76RpeaxqoO6/dLitMgokYQZEH5jpw/VuEYlfNkHchH9BeIoqwvZQBqm3WpLA41cS+K
JnWP6POZCASbzKsn2P7J5UCNk8mtTuXKSu2LOKlGSwszskzRlPtTA6hA4EYlf4eWL4ALIve2xlt1
pQhcRuLPIHeoOZ15AEdm1KGlPkfrIApEtEJViENYLlpzZP3JOrgkTZU01frhoBHb6ftpXUntrkjb
FnfITBNwnysA3A0YPy0KyEaBKwuKtHPGQPh9ufzHT8WjyIB+TnTLycov+7lu57mUnFsp6zJH4//p
dmilTzUpRB9L654QsK8129mt5BObPa18O+XRFRmFyCFzwEX/gpwG0v+1qjpT3zyU4fAqSV0Ptrnp
VYp3FairA+dq2djXXy35EJHiFyXsKme0yOtSqPAITf+1S3rilkeCD/n4+5YHuSrpoZXFJaddXMV6
B97b020ILTVC58GeZ6amfR1iHGF+rupUp/MPoK3Rgm9muPXpTVBYmnhqEgs0uAgiNPIVjFR+ETmi
LuDUSUTIhppewavb1z/Yi7r+SjYeqk4pHPfLJIFh4HCVeZetskhFcln4RY4mkmfJMQqQwFr5GAx8
df5vc7dvY+6PGahffOg2tWNHSIkCrvDuwtRwTicDsbuBaaTiRP0Bf6s8j12bD6EdJvxASPl/oag7
QS7kBV90v9ilhq5lYf6fpa6ooFhxbi/pnR2/pPlHMIFH/6Cp8Mx4EI5yB9up+EsbIkLjEd0Rjdr3
k1eGOKOEPna9N6WIpnos+9u9BmxMKXgi+E6XAj5rn51zDb1QUVZ1qF5KBbsXZW8KVCcST7f2/KNk
DAG6a5LBi/G77KfqUMvYq/J7t5u8R3uosGEG7svuFVxiWuDqdFk40oaaWF5KgtWEGNh6Hj0HE3gd
++o907AvsRK3vxfcybenH+JJeNBNRfRjsV11kOYe5snoHuTgvz9aUSWdmvlcZtfj66BLagAIECzO
r3yuxXtInEZnZxWTPqN8ayNNX25pJ8qtpFb5ohXKMYuOjy8I2MKsMS5RSuO+bQINL0kyNusdbFVk
AV+CCz7x4pD2OJ4EKTEp+vi13zi5ulCIZopM/Aik/f618f2Hgkfppb7+sc9WihGXmnLsUdev24Y1
8YuvJx+CDzc7irUsiOpdZh1r0kr30luIdHxF7GvTdhIJWtoiorPNl9DVLndljMSWv5kV9qLiepch
e3k0DIZu/5JFIfWg4mClvoUDQx7Qk3G15RDHPEe9qzoATxVuqWavodHZpq87kbb+IwtcmpJEYfkc
4lJliojy5nzXSwhIQ5YI9opxUyeQGQpdb8TErK1MZ5fzGbvcKL5CfHiSEEPjydt5vosRA94DfGNf
U2+zBtwgIsUTGDmzuRRQqBdGNHo9xbrq2IWZAexcDuhpE3/wBQqEeSn3l79XTn3pRy4pWZk33t1K
uhOowFDu4oKhlnaKCrFAQ/V3yU3WMAOGzO7CWsq/q1mPNdCNyzIdbGeD/jXusU8Gsp1cZLl9gMOr
2niZf4tcsh1WVmp8yySXyCfcr4c9oTXsHSr0hj1C8sqVXfXqk7UbMOB4etP+KOSwGl6vtmw76+yz
seYZiAWC946+lYa+BYcbZ3RUF6o1w0cRgQXJZAd0zEJOfX/IsqOw0xnqU0B7bmkR3Uppxp3lwkdE
XP0gnubsw5aMLe+QcIHMQCwuhSa4exJqL2Yj3pkdwgpjuI9A8aXAW+GYYQHrqa/UuZ9XKwjCA02B
rSigj2Sdg7LOMreolZAnmi13/iZE9siE3guMNEsxs7TO2OPAJvJ13K3rXBEmmgR3gXZ5fwuTRuLS
C2p5W1hKszLecBrV7aJ7Q6+8CrWFy+d1CRr5LyC7bTB84T6Q7VHUUmyTSNgbuJJfHP3Y+K5kGntA
iXKjDk3u9ZfR2RTLutgaAJK+OXAbVTvFDDL9wigUFDaVyyp+xliRFiHu5wO1ktYLSfJacvsBkBFF
z1FMJ6FqKEeUeNxg6B9tS8SovgyLMTDuN51jAE5gs53cuSknCAV12VIZFGtvRDdof3rQ7GbbQTll
KRBnQKuBol5yYS7fQny0vRrc2ETYe6NjzDFxQ14nLXboUur19DFuEZtnoF2eMdoEodEqVYSLBYLD
jkvLjkVPjVSaIF/wxAcy4p0oemqlEfpT1N9ujeGWWqkSZ0piXaZeU6UetdXOZ3jfmAKLgNIUHLQB
EeyhcxJ2iKaclbJM7MNAbifrRUeltXgWvvJLShFEueQ9FR34WfOuswM9D0Qt4gr30Js11wvHEgVy
9GwjnqkO62HbMCMToetMtlHPYmnhhsTgU0QUEg0AXOOBhqfcfJxZ/Fr8PENNrGABVKaIlQ+k3nYp
kI2k6tj5ZNtQKT6AQBa4vwReOYY59BLPzvFsXDZAcfCXgDBRjxqYwxXPT+8TS4a+X7ovxhm8+2rJ
nScxhJUEvj6EYw+agUNZ81GOsXdO/ST2ym6PkLlc0YPbCp+vbGBFtp+T4Pz/TfsTh4rE6paMFMft
X/FImduul8BaLhuLRCq1+RQhe+CVJPbZ6pmgcYhhPqjLvlgEbHVzWc6URQlWLkttqeJuYRtxDfaC
zALeWPmLj9nIG7vQJjvSXrpqnypjj3Y96NxuzLIxc5fD7t2c58Z5MoDWkHjQUz0Gxi5hX+kdbGsh
bAHbTPNL+iAGIzdcr2MgJpVkaRzkIZeITnI1JzMrf+4LmDn06vhaNoEudlRZZDNopXp+pBjnDbrk
GwN/FjJopbC/NL9u3n1YFVJb8CzdJLp2tUo/BUyV9RMAlfWWLziBx4zqyTz6A1C557XJ/QpYCUwP
Th7tvu4XxmDjZtiD6getdGIXaNvPHd7daUAes1Lznr6TEQNfHdG5Tspv4fIrDIjMlG/I4ZbAD0Oc
QLU8Lhy10HRpLEwpmPIwnYVH5YXEspCqOCvMXfezimaWQEF5/PgVrvgjRmGS0fgV5mkzLQVdv6ek
QuuVMTSe8Q9f6iHcImOH1DaTM7W0s3DKPxwn/lgFv0aZuCtcSoUBWGKfa1ZH+dNOLlnztx1EU8hv
kAlQcqg/DJHwfkUnWs6nZ9r28sJM6RGsT7+eiOOpshTasZMK5XxMn1DpzXJPUOfJNXQ6a/0yORsw
NCSZkzKKh4ZsrVbsTiHuAKRfMWrMvt2UBWC+/Ub4SJW7pm7TUvAhh/9A7CULOW4mwS0ZhcZjJp0Z
F/yoVzyHlJ382J1U3dnul70zbOzQBB8Qv/4jtqRCHBD1YYNAUVNsq7A4Xx3Vnphux5rPkl5oZF1H
Cr56G8+f/WI2r772paZGkjPF5cD9JiENFcuUUAMFAe3jfwH571rjnZFFUtNuuP4oDqZDaahK3LCg
efUs6kRiwLBKS0FIeoS9PYqJUKlG8koLIlnliVbHRV3p4Ag5PL1+pndnmomioTNPsvoMkOTtbqgA
3kc+igchpKN/JBZBu5w1unsGz9vbIVelUqlT72y1wtAwgNkjl3ECOtjSITiodJS+ZpUYIDF+7UVP
1eP59WwxLzLJhsZaWHezyYogq5RfyqPPEsW4z+J1IxTEYBtz0Yr0lC1+u9K96wkq+By0psylplI8
boUAk5L21IgEsJwrVNyuoOKzRbYBxSm/sov3+UnsLwDBIeVQRyNFcoC91VXUoYBDrNclr7a94VGW
y7w9zibFq4cYYAJ/Le/cyWiHM6KvMk2uwEOdZ7Dp8hVFjoqUFxg8tvQ9ZLvJwfmj5rHEBAfqO+ic
glbxchuKg1dW516oGnnLEba7IXGlr3FI0Edokzbd3Q0Fu9RO7cn9gRR8DVCSTAu0bcP15omB8OQu
peOh1JJBnsyTmklgu0IHfcy24c+xBN656+GPVF4xhaccejde5hGu8FkNHsCiL//4O7ijS5rBGg+V
OybEX4qhD7wKBvumkzdmo42uSb4OMIjVNGQ8ZwmR168e9M12wVdAU3i75rRSDtuFZhd8aeoe4l79
hqrg4ICxVGDzJAtGiDxW/XrziuFYNu5iWi9idagK2V5Hrfo1J9zqdP+BSY3p8DXXG3flVn3wMqbW
pmFavGu7XKZsW43IFxZT6leHH3IqlXHWZjLZabvIeLa4as9KqyvwjDrc4BImCg4zpfJoff/sO/ec
V4gLFT+J+AjEjz3G/ekPnZ4g8vTYo6y9IeBBzPNsMg/MnX7Zru+BO4mLUr1qGTll4moWo68p3gBU
JuQye67JM2kOBriUX9I59BNjd6iC0KbD5PO1JnGXampJ61ZHCD22Kd0vfMeMzuzQkmDLE5QiJe53
N5VW6UYfliYdUYnmiwsBX13p/N7pv5CW3hOGd96jRZYAyOdPHQHYy9Qi/6AJkODx5EcO/PGHod1j
0dLSEf/RRgTySjQVSO/olxJNMAtELtMHYMsAZ62kCV3LTDARgCfrQPzBZ8pX1Nxpm1Q5itMZAaM8
HBLlcWZXUjafyIzti4QzoEGFyffK5XjuJbM04XFExG5+/5hEa4zbZlrNKslDxget5ND1R28LfVbI
I/O0QerkiUE9yvF2YDPUOx8sKW36cDV06uoM9WqYSfUlRRpSAwamiTROfiKIgoAHcJ4V6ks2CHac
D2Y9Hx2y56f7Urtx+AuA/oCcrkcIxuZr25YtFdc1b0+j/npmPPe1fmIedr+/LSZDsUo/rsmLIvJ0
FEgrtn3chQZqP7liYZ5QeENV3MhwTmVYhgpL5+g09OeACbKLoW5T7wtjseoOQ7PWDsdlKRu4Aqjv
yAwI77eJNpNGHmoIdzTw20x8syuh0QPYzYb0FR1c/YB0DEkwD1Y6DZZoBCXOdTonRP0WkXZnwUaz
sJW4Ql3cjDV8ICIco+YoA4zt3pBiFa4WBE8mARMDsQqpZiQWPC1LkSOw5ZS7uixEG9LClWc5Ad2G
ROjHgJOsm0J+Xt3mMdr6VFfzzKZ+FMrMZCybzGS3/uyaWrTDoITDrNnzZXwVUjeJHQ302g59LgID
zDGD+RY7ElsuHS5KrAcoFGDkGIlWCyIJEYHawumxlibYWzHEOmPBiPCMuZMs3n92FJJd8wzJn4af
bDTZ8PkAjtLgA+YQLk9ADY//tVyRJ5HV+rNvzXGp+HK00sXnw7kggZ4xWKfTxdSRC+O2Q3Wa12C5
lP+2CKUbzwVOUTV+/rkXAwytcEYbWlVjoj0dXQpDi816kJCihCExNF/Ro/mmJ1THfBCmGxHXnVAb
V5CIG8nUAny+esG3uj/SsFQjjvw7JOhfVSNiMUoHkt0H1U0BlWzV1RyiBTYiIVZYYUPM8PL/gWsT
m8fc8AIM060ihybdytLoYHeFTXPK4KU0bfyRed0rxjUt1IUbO0EAvATdJzRXrx/2yetq4harKxGC
j3SNG5tUPOwpPo0m6yVi0hQV4Yk8qWQRvGMCjVZEavQTd5sNvQwbpPhz8pM6FMv9Mz7+vVPCmjxV
6STwOtFvUdayBeWPcAG+7BcvbRqQnRNF2VyRufvFIon1VyYSlm7LTGlfLcLS//TVkSEZCfwMU97W
qWIErF8NkxWsRCXFQgCHu3EktRwchiOQM2q1wFQy1F0I2LOGpdntG3fU+HZJG4zZcJgV/OsWCvVW
2L+yaJthxcRCFTOxdfszHfAMmr9/vJRTa3wlhUsLmP+rzi1bu0CnYVEr//f0ZJKGv8WftlVLfzzX
hqpuMJC9uQfaFIh/Gj8Vi62eJTFffcbLSlUEujl2XRbMVOxxKdlrYAlsfjVq+j0FBTm1co0t+WMr
oZRj9m7N/ybfjwaXG8rU1bv4RE9jtGuWoB+XZdiiaSXPxO1UlC2Q+EvFo9pOurACY3VUbXxCD3DL
fvXVNlrNgQwRF/sNfS6nq+CLJppoGPXCkOqdd3vypX7RJ2m4ICfyma8fSkkKa4B9+NBKevV4DuUv
KuSvkUuPV8dk1/UnatFvNujTUO+eqsOpUdJz/OrAi50nJ4ufOTQwGXolkGsywhWx3oD9nk+11BG3
m03d6rfooalueOT+no/ztV/Qix0DMcCJD1SshdOK5jh2B9fc6NVEOGC9wQ11h1zVNwJkwCe4zkUM
GcKkW8YHSXv5o+ahai6fgmuk8CgeKkd8R93NwRUhcqSfOFRbvwAuoKyKfNQVFbXblEvYH9qVn/xv
x2uQk6U+OvvAZ2wZFH8FwId2D7CTuhscO+10TVQSUzJ+AMArj5qxf/M1TQQfpPtyPuCWfrwq6ti1
NYVu/9DveMaie3c5SkNKuI8gJNyU0xAYbBmNHZ0S906MqXRT3PuqNHXJReTezTlOMlzDUaELtoUL
LIsi2hlCroYtDSTFJ7mBfNsLOhVsMcoqr7pyYTjnhawQadB27D3jEE06cWVLRYsHxDkCs4Fz91CH
pfzv+Y8KqpuquWq2p5K7+XtZKkr2IRveCtH3Y/9AQqhgMHnYqEOvVgkb2YxwP5JeFliYN3Rbcqwq
NC4Pww/1Y8tyqXRsBhtoHz5Jqg5OXO3JVbpT9Lks/fGn9xnDyoF1xJaJvW56o/xy7d0hvs2IIx3a
U6yWVSJqPgkrojMs/kt3ixjz2LX7ECdNGJVn0CCiCX58+ixXkFFvSkWD/vknCfyOHMCoZv5himPB
a55mot1MO7fGe6WjQwiVpGLFYmkPyFhIBSh2NPQEUNOytCuY2qW91rqr5MCWl2QdUexpNlzzzyI/
XFvKS+VSCIaUwADIBEDY7oNuZYXd2907Ij4J44w8o8HgWRqF9F5zi++oAHV/wApoNXFJDmScuvF0
pGf0nM9LOFj/TRUa4HnDMYd/aSHRYZsvZLdaTbpNGhZBsDcPFsDFWhMh9JIjePoQXHza5ibAd3X9
2JpyWaIhyKrwO92Tx93MQOrGkikBYl4oXPDUTcGBUwHMjVhgbamHDJ01vOPEDnxVHwgzmg7xyM0+
2KQFZi6RbpI6j6GQ6VBNnEzxTA31vEQPb+zCpJNfxThNRtmJBSpSfLqhQAYCF2YAX9BNqqIeczWz
ZWKx7Ti8Y8PT2RbSBD0ifQ/cLhW6SAPIKS6s/978s7gPlVQNZP/QsKjak9EQRJFllli6BVt+MzfA
PnkamKZ/Dh0Bsu55ipdEixYaejRXiMXEGvtNsh9UABEAaAnMMCXqXFMCBQ0G+2p9FlyCWovMONVW
0m342py1DMR4mm/UtId8awnr4OOoYO7C41PmMZUjca+7XhUG4/Lhax3JgRusYtmH7mjkL3JV0sed
mUfXISLSW6+QNQawydntJKcxqz7jeLowq8tnSFyqXpPNVul26wHszzZQMNOdYnf/ez7lppLHKJt4
0jLDY0TYwJ+fBcgOptBJsoDWNYGQH4pWvhHXe7UgM3mBX3PNhYKpkdCe3RnCeN1efNfJMLvEPruS
3WgEU0Fu8mBHKaoB5wS6F7Sj19t+p8HVQk27RqtDC+1lXnyEWjMhSConlu2XR6QTIxKXFBxYI9vW
aE/6kkFH2FtHyaByeq3ujVtcjF5OXjcVBwU6mTZnPZ2oSjliJyP0Hpj9wJMHthgOUbnjN0USk3Ww
gQycuW4XLeeFGHdOdsuASPMGIhsjxh8TVdKgTUaG9ISFPLqshsKP/CJmRVDbH1S7YYmjuHV57EW6
QdAbEDD8s2erguUvmEiZhFiTNfazouIaS9FBUE427DycQqVbPAJwrNfqpLZ9hnpbQcjdxUbJYI0H
l4pGcTeZYyjIoIyxEQR0e07BOtdq/Jji53xVKwfVtl1rYd24TDKa3tdsbUZRvPDp4IhI/gXGA7X5
VS7RvjUaZw/AefUFZnMVSfWh252iOetjYFpO7qLm1MjT7753BTQJJaQ6ky6wtAxsdp2ebSygmtu2
FsryX1e0+WXz4DWsAn4mWJppOKiTo03f+N/feZO+w9pNf++FyP5ejlLlblWKjJ/Rcv/ZqM1HDCAH
Y/Fxru6R2pdHC2XRWR17764F/wOQNgXPUiliRulZhZrHTg2T03nSPrsTpJjnPKYR8koMrqXRbhvP
mRcVqy8M0eZE85ylSTUGhD8bWQWjS+gjgwJqKX/VH+Kb6nXmbI5dddcOaKxnyYjTvSnLlsnuBOzy
24dLIlW/BTgAEFErTfFj8j+FhlVtYsn62zFeyAg+lxV1CsANfu/zwCjl33EtW/4chrKf8oN7AAme
KWYWexeYnopr+kvIP0L4YhLf18v+nqRedD9L0n/inmdybitPXofSKHeww4kAT1BO+WFIICVXEC2m
FO7XCg7hoCB4a/jjE/ZxWHvhMN665bVhn+C4E07Bny6MfWxZ2JPtOQDHcDpSGapnHaLF77ofV4ZI
CJ3d83T5Km8vuRZYMyFmynYi/FbaLPg7TPA/LI5W8fJ/nvTvhWGRjJ1SL/VYwfflqUtHYrvDh05m
pDhWhaNBHCrQKufLOGl5j6gY7vM91ipa97Ds38HToXYucjwwc0UZS3gnwU1zh4iiYmat2k71jGDh
OOYxKjwd+TBD4XUaLEzaKceXK/5C/rh95QaREqivwl92cbJeAyrqw1hqLIhWdTxQGyjrFTHCJ3Dp
Gp0BA9ZYP2Z7Zjdi7Z0eVhbnFoHcFa1AaR8uFTuAVjgw+b7Waq3JUwBe3hfN88niowQhy7SAqGqi
V/tQvSqBoxaUPK01p3tyPRPnsf4/Rt77rneQvT567HBKyRT9IKErYCpS+PZVDaMvk/CbSN3csxrT
qPWQ3q22OO7OG1IlbnCCpcm2kiVjwHwBXOP8mpmm6ZmMT4EAMnZaUqlL3R/TP+eQWWXryIJQAZtM
3TM/qkBeioix8vXjcl6upECbuwqJugxbfAiCl96Plm4fdHqWsVsFcUFgc/CxLaJ1daPgBWLAAqml
lQ8nmwklRr2O6Tp1jE7hxipL8NRAuR/WE+tWY1YH6dY/eD0PevCs6zs+JX6zly/y3al81JI7y7T4
Wo3bPqSwnet0yARTbMiyrNudWyH7FC96UhRMWxY54nI+XxPB6ZWCzu687jq/6+oDjX2bj5X2IQ8V
EJiL5CdTbIFSFvJ67gcoIxi5xIAc56ly4d12x6WnvuAXIifc7CEmY7REIlkoNE6uI8Cq+ETr82Ox
qwFblCI6FVMaZwKGTHovzbwMqeOpi/yrKKapRZVFBHcoCoWijswRHB7OtqbiWRHnMTJ3FoIUNbM5
HFh/PUEyyi3WBXYVM5kijw23fX+5UVt2h6dHnn84S/CoDAeKqPcvgor20fCkuxIlx1mvY38MA/Z7
tVtbKsr2DmOiJTVMT0WgWplW43Dxs+NXPxPbQ1SISibK4WlT4Nqb1D0FmcLd8PJUI/paZpCUucqE
6n2YX1TmXr6UJgo+cuaAHFw18Ms5oMFXHr0RxjEcmcgihHqVx7mHQZqLYwBFR5B5DVaP1EMOJt7F
DuEX9F39tWqqNnOu83mWAhQeu14Xosv+S7mNbj3xGL4m1EWkv7R/tLyHdXxsc5ujQS1WG8jcwIZ1
NWS/rDGdHAa5oqzv4HHAe0RIdwgJQ1FS/4BBmwTWdWXPVd66qwwQcPz9/k2NYVkO66kj3LOfMGXn
S/orXMAnfKKh9vo3nrLg/EXmcB92vNJrejtLE6vPyhAVd+X39G4G1viAC4G2RU2JDnnsnVDyoAd/
byC/TNu/o1hjrsjggtod1XAYORQjGY0W6oQrFXA+ANnEAdoReACxImUwrClzaq0NcHauKL4/mPLV
qN0dG9TkpPwi89XUTDbT2XZDiCPTx9a0WcjplvaqD3fcgFx+L/60vvcRDq5DbvysIPRiog8KJ/Uq
8cd7RColLmv8dzoL+xclNv3kyy8BVDF7tW9x1C+FhytMK/6j+o7sMy4j5FzOg//+dNLkHGtxRXv+
UY9U8YvuekX94LF2miLSys8Ug5t34vbZ/PPWgvlXhF/5KVayDSb4juSx4s+WK7KcGYdFdkKvtYFp
i8V22/jepC+yOQxlKLAmME8oa8nm1+zrBWlLZtwcD7wTFyEBqEkX/217j79FpDHypkYuDHFh/ryA
92FHsDCT4gEaVzxu/1iJjlu6dd30Za8+Rffaey0LDAuu0EPZvwz4wh3xy2epWszPzSesGipn1PbK
IwzlvVm3Qj1VYqs7cvYRhfljUvoh5EPOLTDyLDluogy4UhSu5b97dygOV1YZ7Q3TO54d84nbv0Mm
ac9vIu79+N1xsyCX89RXoyHnUlN+0qeIbTLu8+ViezDei9P476zj7FL4ueMmj2LTZ/bXW2voYn79
SBSEcIaUuaoCVdRqyRLxJxSnFqQuuVrWXorj/smjiuaeHaI/BipdB27wV8LViKLxhuKlGu+/Hlec
GDhLgrp3kRqOrH4a0S+2R7m3W0hlUt8vEDCdUDja2EmeO/Ku/TJd7k9QydEib043fTut9dc0HxAT
Xk31RcFKB3avo0f/tKMLDY/zRoppzFjva1yy2l1sZcM4jEnmsjuP1fK+RKm+jxuPDqRv6gyCdLsb
Zlzy3fEQQMJ+ZGRFRdpLuVmk5cqZ23AgMIf6qvJHWXbNHWEGerQLd72rhA4EvuvkeTMb2dgiSmct
0Ro5afgicX3a1XXZaT521tNLI6xyelcaNpy8AVrFa3XTPHnuRhqWWG+ME8BpYy63CZLw+LoMzfoZ
Uc/4K1E2GMeJ5At+05a0v6rkhKvEWRBRQbkFkmD8IaaszPH6M9zrolCrGQzKpuyoV6HkThWT2LEJ
UiUkgmBB7+k1jIiAzhLeb+LIGsfMXchjnQRirnwM2w7WxQy8Clyb6Jxj1aZp1HXW0XW4Ar6wrNW6
f8bCfhixZHLL7C6d3v94rRkO3J4VQwDmFNcE+8xNR1yeJCWFqPG37OiQx1NaHKY3Geoh8r4L2REi
7+suzedvZkEKSMOJa/jToNmcmNo4QsUfhvUNB999Sip+NNMCZqaKkLPPuF4W2c7k/7cml9iOoDCF
TUxftOXUk9dU6LLW1GIQlVlBzw5OsKjh/IbHM8Oh1/hVcZwg+NRYQ3UNF9k3EBmxy3KDF+kk3F3+
3cnH5R9tDpUx3m5LzZEYqz+7WQsFFb+9Yp8zdQTIkygeRmvIvk6vt3i3zu7ToRBSQG7g+w4Kpf3o
H3Ewx+3t0ANTEEvbbWv63k+XVISl3T6sJfGa+RRiJpEYUWno8pPT1TGeyCLrQLFrrYHjAfqrX0fm
BeXOhvtgRyj0dWVWXDyd90BlhM5VVrEtbyMUghsRWDEoEFoO+K7JSdcyphDYvVkwB33QPlpiB+yp
kwFbplCmOtkUA/B0NjYI6Q1Ta/4t1XPM6HDtoGFDGBFaqwoXigSor2NFZYCDntQ1lEX4xz4ivXK1
76mZQohYH5k4yE4gWO0mp1JCACMIiu6eC+WQpGvAtuhsp3d5GY45Fpe46XAWxc5yWckyf5vl6ihK
8TbNehA6afJUKq0Rgo1Vrp3AOgsPgpjI9i2VpNFCPSdU85e31cgpgSP3t6U0hlz1/58F4WgVfdO4
E26sP9Rn/kdxsZXQPkqIBYXzzGIVprfnnKaQWe1ZxP4g83P0YTB01PjVvggmef4ObRhSOc8d6WeC
vFPPsjvgA/i3THGsT4uQISqYSbQbDu+iluHYO+fI3oNULwj7z7Zh0KCJcUnE6G5SmRCNitVp5gG0
on882I4VU8v1qWPUMnvZVTVIED0lD4e9Q84J0aWmY76JixrLXNcCXbzInlP39FhScZg7jKHgdbc1
jbw53hWInJ5OPOOMOCEPxSoSmiyn8AoYW6dHq6Xlgsw0yuUqspOSXeS7sAHWDD7gCDJR77q0E0Oo
1lazaJlrvt1pgbd2RGCto5ELZf1wGB/HOvrUHK8h41jAkPx0U3BA5gyCS2r+27KoD12ydm1Dr5KA
vBMAwb+gfbtE6nq5SAmGAYliNb6G/RaquciNwkkgh2Eq2cR/PPZ1sNRRAPtrPgk9tuOKrgxut6nN
VLRWluOqba9jE+34IPF6Ttk+BKk9GSAb45pVhdmdNLzJq2x8ybi2xFG5kWVUZsskF1rKzKqqerlf
qTBBttXkgPlfsiTfX+oY9WUfXD/98xkBkekUN5uaotV5b0+w8ebvNlvuoRYexvdne0pSjiihPI8I
iDfB2W85g5AY/rAhcip65TyqvxGnEtL/MzyySfols5NioDl4sIejo81poKGx/ij+mWz94oU1rc9M
SM/mR+85LFkSjA80TARb/eAEGhqgFi82cT3CWENUD62BhMvFtCoVckLN9WDPVFHhP4Q5n0FYtWFR
+LNSt+mbt2kZUPdbzNlJab7uxw1iPzaoAAai5PxBrlus8hVlgIdTlRJFlM5xgO2iTYvb81OfNZd4
18yMQPoQISGHTPgeJ7guKav/0Qfo6lGuIfdGS1jWG9DB/0Qj2p2K6zsHpowHOM75KgAc/yXlvb2z
a6FGKgF2mQ3Yp9u8gxBtTX5cK7THOqzC+WNIEiAvpHJvBat56ceh9nfS6GtJyM7vTaYuvxs3VdPW
TvGYildMI/CVxCmJeBIMQMS+lg2iwcTfTv/l8Ml3dC1A1fJeQ10ba/TKlaFMinllT1+mY57mSpZk
HyIwUU/O9TQBzlTDlacqPGfc7iKa+/EJvNUlMiRp/x1qF8Y8laqyJj/5qicE9t7cSfQxoPMUYpuf
aCa+yu4smQJ1busiMVEI6n1cFTo6+heEVcNYAlgYwktSHYnZcu7vSUsQWgeZOtYH16HSItTY9sOq
o7tQ1VaAGc4G+06bMJ930Emb7+j0W7mGSc4jpo38o0A6rj/dabI36h7vL2sa0mFF85MsWiPe2eAd
mrjySv+dyjjKcO29cza1xHuc86w9vcJeQ9fSXnGjgfTRqFd/6bA58ZxG2Pfhdmo4selMcnLDMAye
AWx3tK+Q9KWpNKEBmqcywE3EVydsYq9Nw2PRigy7vInxIwMQ+C4StLvKzz2EGTgmqBCu+OR+ZbFm
Sly5pVNxpzGgl4ISP6ubw+oYXXgSCU7GcTCSsXdaKR29RaUJLWdWIxPZXcrMlq/TDCNF66pQkG1D
OL8H3WD9zSHS2z/m+asNwHO6BPAqU/EJdN8oEIm5zqiyvxx9zfkKXjvDYKfo6z5426+lO7t+tcdx
ToKtko33GUnrP5DVjapJhCAEUWbnur62utNo+l6HvA5CVN90jEwm6T/IJMoTXtbghiamWckypR4E
5gLSnJ+PvyBuE/dW9hMwCNTNpLtkX1UqGPNhdVwk0BcsMNCvz3iMTokCI4plNE2xJiukVKs3C3rV
OTLDT2dof13tqSPI4BA0nGISN+MH4y9CkPXViNR3ykVpJv8C3eyCuvbHF3VXt67G+vlNIouzjHeS
H0yG1Zm/kiSZLwPGQL7VIxGBjzsWxljt/fktxbJJQWqfugkls8Q8Dt3fy+Wywh9bsyV5bHd05YVF
5/zbHgfZXEXlHOl/4Vyaew4hKcUzfW6Skrot/hLD+MUXxpRG3h7A/+BAndRVaPULFADmCrDl9lF4
X228pT80yvm2H543liBegExd+rNs/XColn6uzSffPicXEE94zxYUUdo3703wRQOAa9pzXpmtNP1A
WCy6HOwKf2UZwUnmMvcM57eN9oKyvBKoW5jv+EDSQ0lZwDOhyCFW3hX1hxYK9+yFJZZjmet2+n6E
1dC4c4XofBDTEZkS/EZnKJg6qwxVi6IOQBesm9B1VQITqa3FYS/RFdyinm5LhssEiAO0IVuHtuSf
nQvD/HCWll+SAuie6me4NJbmeEaGzAiqGVWOb+L53bIez+/bev40VaEZrr2DrKpdP85hElp3DKRE
2vY4vgLvrzjPxfd2+PAXtaoj8DCoHF/iR2/j146I1ysPP302J1Z/TiRkzdi452nGCl6Ngv43bqnz
gJfIUCZW/y1F68MhP/WeCLZgwgPCe+x5PPTmMbz10vkCa5qIWER8Wa5NqTHTZDwcRxz12CzSrFhW
hmAwSEzlN/q6Ugl7A/u9SwRTG463ghfyqvF0Qv8XVVPr6AKfJZcMnNOErBPmcZrU2wn6xy4Ih2Cu
Dw8DvfVKkT8g0xVc5tL+FC0AKmoI7RUui++MCZZZ0kuFttT2wGY+Ht8SkDCIrO+wC0c3C/5bYDaJ
3S1+3yGUI8psT0E1TvROEUeDqmNVJlnmtAbjJbft59iN1fn6sSPfcaiNtbZMZIm6/D79jUWYnsg7
6ylHLw6uO8x7j2nKHZriPaBOM3/sbtukfk+v4Ei50KpMj5gON3PIk2xTD2j+2/pG1OS1/W9i8W3Z
UTOCgm0SbMWYl+keNIzKNA2aPQSK9qA22im2hS9xO+bF/O8WX1dyYJCTw/QQhqcS1JzPMjFX0ht+
AJjBL3/PBTPNYwQxOK5pKdILqoNzA69gxRLXA54QRILFFiVU17DYAxiHynVqk232SwG0WTgPOM8W
95x3pilvH3WEVsI9i713pFPE9etGC+qgc8vyTcxk7IJcxg9rl9abBZ1Sgn/CsiQ6iRgCh1u88MMx
kiNIEPPjJdJamTc1JDUYYYxaVkyFKmuLHko/6bl05uBxHwmpDBvRhG3cIVtuemsAUErb61ic7zhU
FFyo98L9D8AobRnnrwx+QToW4Kpnpti4G1fG9tmP3MferGI/iCEnZOJOkpvkhTGC12YG5tIkR+vB
FIA7+3JpRhCkZ+vbhcqHMy3CausEapAua2ePS13SWNRCHOXqQqHIlorS9HM6mKjc4HOYx/+Unmeh
Li/N/yKDl3kBpq7HmMbOBDDqYJuqh+hN4DYGY0dWREeYnAcXSzwi9DQGcvdwWsNr7/u0D11igUP2
EGRfJa8K6rWjgQCUKOzC3PofwvulOy4S4Ps4vSp4Cdg1SeNXSGElI2BnWRuwP+bpNWZcgzPLeZXW
VvbspA84LWhM3f0Q1KIN2q5FFEzyNyJcecLN2GUYAep+qtciRKWEvj58LMmhmlw53382wc+UfvgI
6t2nBUw/4LrufszRet9CsQWZDlMt4i77uqSjRwbErTSc/JUPsTRzaL01oGpG1s+K1Ukwvt297m2P
NSFmUa4QHdP4BuGpL/APFZ1RM6qFMkvO2RFIQnCgsqXH5giVaQdoT2jtLBuULUdjg5+qu1z7EysZ
pXk+hSWihr0l+MN4OtH2runeUF4YJZELOxNNAD7Il57g9156j+7PQxTLnFa2XVUJRe+iPM32MT4m
IOWxhCMrJpRIHb/u0G0ii7MpJKPxBUc18eT6B/1VUjQQhAE7GWx9K1H/xUG6miqjJI0wOhHZ7XVx
yrgPFrG+evhO0m4dertHQjXqbpPcksxiKkM6AKGtkpqlqawm4swj3KuPccaciaH0ttjXnExb2xSA
tUtk9TbDPxz3FqtBxU8rQSZBuvFwazJ+dT66nJ/jAgVtUS0PvbCXOEXy8bn8s9EsvRwpDq/ibRbV
x6P9YVEqS0M7vgpi4HSKECgojROr9qrNDuXA4nBbpLIXBpIRwdo05hfJlgX6geYg/JnfX7AfNbUa
M+/ZorKuU8nfMkb/j7KTk5iDaCAOnlPNdFWuUTc5cwwkIGfyj/J8/gMYz5NjCNMHjzUiEButLuX7
7mymzVItZ1QI2JY+CHcPojpiFdsIiST2QXg1ab1E49wXAckAnLg/KC6B2IU5vllYaZp9aoxnufPP
EL5WW9N1WTQofFQYPhF5ECFblwYRx6FELI7tXBZ8s3QygFOZwcsbl5LSwKFH/fvG6QTzpnNACxR6
bYgT6dtQx3xVbhQ2Uzu4iZ4bEt2GooM7MlZOvduIl0/b4RFYmvxt/MGZO9K3Ig1dc+xHDeOZORji
bWQvWqwQawp/dSdvJYNf6nLcZOGuVgUbKjibVNTrer5v6FId4KJFJ4P3Y7orWCfhlESctW5ZxFK2
Spbq+wMkT8sWHhdLIVakHAfoXSuecnkAs1txvs3nfbln/g1sOWP8MyQiT8XTSGwBUziyFdXkxYHw
NAJzpVBHX0U3IlHtBPsiH3VBWbhyauXo/eoic/anMnDheW71VAUdInkQZkmOWUWrj5xq5iFDJfX4
LJrMpTpUm+Bg6iTrv3fC4NYeQF9iGamgJZ4UAg99tgnBJ7H567fCO9AetHofW0WUkCCSd9dvx2Rb
zrm+e3rY6O2GWXPTHyyvme+6wSV/ill3iVQ7NFb5xhX2YvG/4Flq/oBxjHD748qBj+c7qN9yJt/Q
67R4Uv/J1dHocRAvK7KnrGtTBtnNvgU+N7TYQXwL5rlCJ17M9l/st3nEm1igRyjkRloU7RsV9G3/
5ZVzxhgBHJQD9PM/RJNmyKzTTVadrIEzlPT+DWZDOnG0v6Drrr9w5k2gsTkuxqc5alvenYrGmIAj
AfDThtseeUZTAmy4EdL2X2gyI/FM7PIzuY5YEHbVZ3KbbZ5qvk7nfSSbdBtvRSQSt5Ub+ffB7BGD
U1INR90a7UHRDmBVAihSMu9+OXj6zOhlv4TNRj0TVkaFqu2fOujAYQoOhrTOYrAmj8igir/MX9aK
xqh6MmgxB6wxheF7yx1hprn4WKV16qd81CgnNxGNUlaWbNkpeQLBYU5JUL+sIwKnK6vMCa2DUFtQ
Wp5gIVXTwtH98CR0O55Kg+LQCjMCgXEHkCKqzfL1UwOuWzSEyHIV/hxVWQJa62oxf5+TTlikIx/w
t1a6s9udWg+26Ar0NIA2g7sGF/ySZj7zoiPFChYDCPv2D43cCmCRgKxoax1M+kyWYVrBOf2fFNBN
1QBFxhtqU0JSVhgKMVRYg+Teg5MrrNceawL/EFCI9LJBfF1Zs4fcaPEP9GHqMFhM/evYAEpRkTA8
bbbcBQlZyZQqF1IQw5djiyECzkOIdnywbUh8qjBHfkacHjp8az1xH6BS1oAw3wd5xf6M+ZEzzwuh
SZU0DnEVXWSVxe6N8nHfiJqrhzkJXOpAsPHROLbkYfpbbrNPPcZwtckJvkUu5l06alQsOiHN/x47
3lFNSA3bGfr2YR+6YJBA6VuaDS7yJMvTXKRuvp7tkHl8u0KE91ZWwzRwQPPwV3Tb+raoYgw7peKM
yfTqbd3N/4rly0jexvbV25G9RhS1aoCUPlUB2L/N4P4USLEZNO6AkqZBx6CB2RMzBH3AYBk07Y6D
TqFQnlz1W47uTlmNqsBGb6q4H0x4d+g6YDrEt4oG/7TWFiuguDLuRf6w1XCy9d7uLS3/enlWUuB4
XjEQbGgGpYFJlOBz5SfwZjpYMbSRBcc2Cr13krJNjkTgDA7Tk4ufPjic588fv0H5vq+oxD5QutjG
jvbZQYB9nNVN2tIL+Fxfj6i5yYrn1TTNH7Nc83huGb7lKHqeTvCwovLmrrJMw5O+ba3v4WY7xc07
tYYqi3fxWpYf9SYZ87OC/VgCxXNQocWwkHjnuv9Of6LkKDz1Re0d3PnCx1mKJabrNyXxa4+a9DKm
N0IZWvp2RXqQ0H39MP+4/O4kyBlZJ7cOHjjReO0S/CS/oeBisDRu00JD0eITZbJ4jZ89PYVyBymL
eMfx9J5ZUlMrkGiPd/U1PO591uLsUJ8eEx1eqcUWXw3i7ywLTvNbf1ErLoVJ60nkQMecbaAfOkIx
5ybrrSmKkA29HbqmQ3zpZgcDjKHeg4PZxoqbC0T1DzJxUgOSvAogBEru+vGjshUMSQondiY9fl2B
PqC7FoHe0lR04M0U2kT+Gpm4IJYQeRl7WXX9VVz33C0f1hjO4puvksMAXc1yd5lqAFfZGTRFVixO
2FkdIrrxccPRU4nhAKdH1j3weWDD42JeyazAxTR0PCNRAA6kb6oYT7XChyTHm9h+FXNF8X7A/2rb
xBnODzQWn4Shjm0jPjPtnJ/Xke8965xIfpP+Cl0A4brID4SwZ1EBJb6WS7smCE4qC0u6MHZlT7ry
BcAfZoX/OFmIdWBrMFufW9vj2A/1MRe1jdlHlAZhLxIbqPQd1q8srK0GCUb7JINUWbyL9aDqXIZO
/a1cM3mEbbGsiJyp4CKWvJO8E/NlPDpTH5xtWuB/fapZXXBeBr8/S1f/77+270GMSVEFxHuZvy/J
oMcfGdp4QDYRTlVmB1rZhJxtYCwfbjfujn1gpgotP8+k/2COyzMJ6YC1nTa1bnWTyGSFMBr3VeHn
jZMLQKZSpfWYJ8h+13ib8QjfEXFGpzvDuUd2DTCETswhByk5NuQw5yUDHvhfkvo6SPZdF58qPWYv
ZHnthsH+TyprJ0OX0i/JmqZnv6TMf/5A0eLa6/eSKS4pAaWOTDS65deW4MXJzywYL0Y/FojX4eVP
HV/OJv1dra5sdhBXInFr+Lj3uROjUIRJwYtCI2ECxeoo4Ljv4ky8xnCqVJzPH82TGSrZ85V7kD8x
L1Om7qBnHTjIe+etxZRIXBSm1EmTIbrtMUSU6UyoVsTyPQgoz2gt6PWKR9q9ZYRZhAgahiZ+a+D9
BWRD1rQf2iwBqcC4WWVUhJIjuGIxHbZhlCp6FX6J0o1uJwKCT/rNwksMZifpHPwKu6Jqt0YdvEsS
jxwAPNQuSR7bLkzJl7578YsHSlvsKQE98itD2n1dm8uUwpCT+buWvV42c95PjaKzNAQnTI+GreOA
VXZL6SSj2razgRUxqK7quup1O5ZmRUFXi9LQqvexLd3E9x483ERRG3ah0nmCOOT5WnYxi9Jk2Ixe
+1VdOEWK6X97fsZH8JSCKFyAkYsB/xvN40dyrvswRzZquGEzSrm7f4VVSgepQITH9LYnM/k+X07y
SYH4i0BPYmRLH9YW+WajQJFJrca3txE3+go+ku5aoj2RZ6X+wv3wdzxqRiYomgKylMTsryO1y1eU
4B/DxQJCc7/IpNVpQwaxa8yIxPv/WXxAH65xxqxdb6kweI9lTJDbeGJMizTki3Qj+l7RpPnC+oKR
3Pjhd3Lp6z6w+J5pGn1hWbOXHQQXlmFZX0srq+kULoJMvtLSmM6cUlSVUDZNGXMLzgssI7rTbPZ1
0eVC6ORhS8w36pvkHMRBNAUSN2DXBWkYhCKYJblqfzhp/2oNo1usyRIpbTt1b3ZJBZ6Y6Hd/uGaJ
auapotOg0MTjRed7Us6me1Qt2CdxjHzZoMr0OT7QmxBTupPQJ8J4E2whpDNANf3DqaXQ32YSFDkJ
TDG4+HiJoMjzmot56HFKCSmgXCc4Gn/I4eoUvNzwYF6J1C0t205xuooYTdT2pFm+Tssg8NcKJ2g9
yYUTUkRT6IxhGu+SDGFfvz+dergezJXu9M1cl7ldB1FXKnVmmWxJ5qY76tO9CNTYSoeErWcJtjpd
Apja9jrX8ONgrwsMg/KtdyHcgNI5oc7jcoaozNcEocmDuAfsHXUJ0lNBMYxMP9d+msLtGzAwY4/r
vbm3Huyw1v7HTQbDAiX7t733W9osydI5dA+adWL7e15lPRqPUEoWZwXD7JFaoyS9cTBiwQLI7qoc
HIhl23i/48oddL03rqXFUF8aQ0Y8DuxYgmNn2n+K7qNn9PMHZhPPyrV+8Afu5N0q63tk3fNUJJcB
7cbbq4w6ky6n9wMLB+b5ZSWWUgCdDoXkaXJ9Rg2jtgTAH7d5ZsBS2LOSp1JtTKfQ0YqZTDL+gUq8
rAtn58fZQiP08yMJa8IjL00MlNIDgJLxuora0JzM59Mabg/mvYG7J1bLIeK8hkGHDe1jpwyYpFIY
0A/0YdbtmizSbQMOekw6NX1enEAQbb0Prapu/NyobTUzyDeqNt36cn9arCGy6gV9wj+QR/+chjqU
o0ndFvXBq0ut6W/1qcj/Mlq24uDAwyylaXZ+Jh//UQe5EYkqG1CZzOnSkMY4gGKe6T27mDfXGAsc
G1VAGgkDKOVQyJ1dQnWDiVxGyoaZvhbLfs9oM8Klvt9eCExJf6mItMK1AjgwsxpIUHNJ4ae9vYVh
nODvcV7mxKK9ZfSjJAbb2Yi2jDigXmEmon08MWWeooe1ploCsPAvrnaJIrKwVOfl7tTj8TrMRM6s
/i1/KtnXK9c9BAhyRSfQxMlW+UHtswJqhjW7Pxv7NqKCMC1q44EJn3rVZP1kMrBZ7AOnkdX3hOX/
mN+81QZ2XMEIb95lxZbwX/ZNZXEA7VIu4kkSyj7vKxcqWfEUXPi7wRYNhA8bOsGGnDNNLCKV33gl
P4mGIB09TD6DsSeQRpQSzBtugUCWN8xlrD2T++whhgibXSv+76a7or6uOOko6444WZCA19pPk7k3
UZ1zbFq6DHdQ9HWQ8/3E+6mRRdDb+9DSv7ehqbH02KLQFQUHElTnO+vTtGO/fQQgA7btoUkoxfdp
qbcFirT/5rHf8z7BKoAFIpZLqOSXyi6ZBSy1+h+9dC8caV/44NfiwvHMQFbQxda9oGj9WJP9kNaO
71aBhRFc9E0dXH1XXXclh4+I3qGHbwG5ijx9KIkuylOr4UHHQOatYyKGU6ht51x+2kdwJpIO1Vv3
7ih1C52bY+74p2t7K1YN3XabT+ZrAdpT+Ybug4bjTislDOtnKK8H6Yxfmu7Fy3pQDqV+qtJW70u3
YXnlwwPo/6IU3sczrwDyxrJ1oVN4YuCQH6tk4UJ8cMy/DsV463mu+TRsvfqbgRnxnwXpg7Hu6WaR
Br1ho8jTIwo7L/r7yH4kcRmzevePLmneV9oKmYDCESP5RtxKSKNhcKMcvhkRwfENO7SowawQkX2B
FwsoKlfzg6i3pAFzdRrgh1ul7lDvnU0AjAI2jcCizG9Xs/y6f7DIy+/BTH0ZccUAP95k7m5GKi0h
cvOwTVpePhNwk+5NFybDoPvyxQxiuYjn9YmSMSPxMclbjYzpQncXNO6pOw8PLa9brdqtr3E4L3I/
hqEXIo8on9BDhflL2BlLwu0KeyuE7thlsAf97Woahoht4Ir0Acq3vnnYcDUa4cnyZKVCVsNZTMXK
1jkBFrmynQcMdhMbYcamlF1GKN/T5LzJ/EF/ICtmY8El26kD4rvrgZJrW7qwjup6LLqLzo3npiLu
0xJw76qb9nIrmk985J4/pGnfWXGvoZycKDVbohGKjXM0lgtCXfbmc6dxYa/OYDjNbdtXuVM9O+nD
xVWeMjCBlASEyVydDxOrt6NpC+vqLcDX6sqHk38A5gaBrzus2is/CrZoolDl/xDLuNqP7ebexBlo
uUmoqpLrDguRAoZjsmAxr4PEyil6U0PA/kr2HSCQxDXROAqFbrRuuHTN9AXY+XqSVcKsXKPxbLzz
dTwHwOvKnQdViiMi6LTaNN9+Rxy5IGGcwRAGyJ863IY8P92TKJMO8qZ4OLDo87DkZMBItTEhboVY
ojFrNGqJ3+XstTlp1kMyKs6JzinpFthw1zw4joNOATmKO1UzAtU1OcGJUa4B8qxoGUlDaTw7l6DT
K0LrJX8kayfxIBYPhIc0B1mEe92cJ2I2ifSHKsGbqO03FvjAdoZW/7NelBqtlX8fWpc9MdfiqSWT
sdv+pCM15eSB0qwM+wNhZMUJmuBVCuS28Eq/ETz6vkcXw6APHE1uVsau8Qbp8piy2/Ex0/PC5+wJ
p49Kxsfvu3+kw+yrKW4McUyjChlRtdB7kM7SODfXjzULw0BUDcM1zmRvlY49FITw5sB9CluMoQEZ
34buAiunSK+CkKiSY3osF3mmttqb5n56caM9li82Mw4tfcWgcvs7jaDjaCJkCyMPUU9Cs+qiiGKV
ryNW4UehxySlGgMIN7SyRmnIwF70ZnGdFAMXw5yedLF6XUiAU+86HLVsY6tFNGw9GUyTR2lWsbLQ
yv/RbXve7Kz7FBctFQVItAERG6XCBS83JgSLvB9yxcX3gVJnT4YkYJ5/hj++D2jui/JX3M4NJxmG
3m+Mt9Tg3tthnkN5BDNQDE4Bq9UYcCKfHkU4hYroJZh81EcnvD6GpzLG+AYXXEj2vG+vpk7P1xoi
BCNKYYiATxnAhbiGjGZ/XKwKGMaYY9S5ZL830bxnulaKcYO0O5zVdDGEnNx5sdF+YKWI6uesve0f
9F6S+mxU0cLfYrTwvyS/ka+MvKpSwWOMp8EJ3O3btMbYxFdyO2FgynYR/W8kSGypKZg9u3oKUh1/
dVdQM8FymwFAueAQGR8krpevooa//kAFEGS4Cgq7yQGiw8ZIa4ULlbR/0ilkV+i6b5gfFRrFW6cB
SO0U40907MDh2MlZinfD9gEpY2BPYLv6sIxFglmjdGndiP1M7STSpMvmod793Ytq/pcAJCb4Qi+u
N3e1P0MDnMp7SrrR5mEqffmDFrzwSzPU/9B5lrIOkDMkRP/BzGjcVosaVLU2MH6x7SYiZFGQaKoX
fV7SxLJUSLopI4hjSSg/jRpzu/Zk0yMx8O5RK9tkrFPdmwwpBL5s6IzDxBHhZ3ArEJdAhc8+1Yyu
EPE80MTfAQvy4PEG4clI3ezLyQdCFCM6T21D8YL2wcHmh7wXh6hoJXyudfo3dSa8aqcB/xhYTjzL
E6MDReeBhEYppj3rk9R6ybkcmSjy9IPG808urD4sJfaDcJ1/i7C1dDA5NziDrAEtPcubnzAfuXAm
vrA7wtmsO+xe2MnUj66rN8R+gHwlJCz2hPt24OCW7/LGUi2oEAOlIc7nu8E4AffvWFS9vrzvMX6y
pQqVA5pQgyjMtI2/RiNrNEwM1qUvqN/+b670BrDFfmiwrbtuGLh9PoXqrnGAXuykXZBd4ivND+di
mOWXgtBWADy+s9Kjrs+c23WvRwEepL6OnYrMtfLuYT3uKYqhRWstu8KfZrXRmruIg/8lIrSV2Aoy
jw9ju277T0gZ2hrTOx/+piJASF1ZKdD/t+mRZsB0WYP6Ie/21KW/Ns9vuD2bfgr2tcj6URh6j5fZ
kpwnKxoJEhGy4Ei8E0tCkCthmy1NPnYXuAI5uLI6HEqFvYY464ePsFHFB1var+nerQ3K/OET9OHY
mXQBKFLRa2W5Y8lF+onTVddaN6Dfz7IngQGW1Oe/d4Z0mcpctoZsVtb1Q71T1zuglzja+Gg+uQwX
GZ640FRJUZtUVSznN/NDYi1EQ/rxO/l6tAUFnLRLJIRKx0oxZO3jsFmfm0uuXVrUgnGFOLWo7yDE
jb44l5qaBw1rqKCc6/ter9VZI5UG7zXmMa+972RzCWCpyFKQRRBZPyCBleqnUHtB3twoJ2oi//Mw
KrY4zFYyypHB1tHHXa/UCTjVkK1EhEKkZWZbgRtKcI5LW9Zki9qzMfUBxIMVw+eS7zeKEUls8BXp
urJ/JZMxX4H5QS71ud/RkV/RFUuwrJxYqfsif2Eh3yTVc5uLsg/FPNbWJtQiseDK/pVPzj6dNGBa
/W5Sv1G5zYOk9DV4VqVJORNBNbV+IlQpSxhnXYsqScHF88xK7gfgxuRRI+q7pkNE2y7KqGiJ+1m8
xN5//ZD8l7LpbM+WyRn8sfVFEpcjSkbzbcW2BKQDIqzFUA/xgtWc3rrATMRbs8lDO+NTmQeUSVjD
duwwWQyoewwBTPbLUAgm06DYpi7A84wwyIsbYYMI2cHqCiKjzsJLgybl9BXBkEGJFeEE5EHmuK1+
jqBJYeCqwsuISuf9K5/4T+zY026z5WpCA9bpd0D8AAhWS3hFUTPEWP9EEcI45zCyXECJ/sGi2L0b
M2k0gY56TgH9hH0bNTsltY+WzRgYAlb7Q8BhMuPl2/2y3ECX58zc/t/zsJ6paixLCAL1ZD3DTt+Z
wk+3zwKzpHaTLEze82pJEZjdVDle97mQ9uLjRxbIgJBk5JsDI6lhuzeZOaiOIhUQc9d/Z4/eX/v0
Uzrdc3i/5p8X/WDBCcS9jeY8TSt5WdZjH/qjUYpNi2ZcBEjKDpHFch1vYBTFRM8L5rkSXSFDJwr1
4oTKy2nLmj71I0+g/wRlfwO6iv3xaiXatNrv2KZRDWiOG5bNOeWEP3/VrfZ6MZB7tSszrIpYvSK3
4UjYAMMZ02rZvPCl3Gn6TxVb8NM7uE9QZvmtAp2U5uOoxS9tYG3ZdZv4TLMe+egY21E6i2SqWnl2
V7Klm4RI6igmPII8C23tOEgf3b5vOUUmZkDHCXflC8TxGDxdcj1S3tiULX/KFeAdrvXahxEsDflN
9Y1wtp27/ARHzyfw9GDcTu8tbSeQLx2BilwcpsmANmTSlIoS2AlrfFxcFRbD0llLvTDcAV3qXcAQ
eT6W3AWG52F3FYK+Fg/L+58Ku5Bsw7tLfEWsnI58PedCNGimtKs5+MsL7DOIVzMWghIumWkwRRtH
rEGr4B8hsJlHib02EFKgonsTY9JyoldBPUHdLqF+appWlSTyTYy1uEZ04q1NUwRTXpBRCvP02U3E
bItoTZFD4m7fRA501st4k0CB0ZcyDaMerItSLdLDvzNGYdzHsMmj5dIOPuDKYt9nGxTyHS8ZS+un
68IS9tWKuD+P1ngccM4y9EoF97VjoatJ2rQpc1wz7wQOYn3wRmQUQr7AhQvLZzZX3nP8O7ds8LP8
iGjGxYhnHXjm2oDXSd+e2S0TIDQaDbV+TeZhUAGc/dtHSznd8vnhDjIOiPF7CcOdNqX7uHOwunyY
6dB1pUdXFibdCEqrl5hYzbHwUVmc/UvfIdfTD2FdgdLmPuPI1bo+7zoNo5VQK66rlQOkUUKVbA/i
KVJLjCQ1FnDulgWbIN1BB1gFokr7ZLGm6WV2vPdp9RXWDvkeEeWbhTtgjQzGHW2Vo5PrwFrdxh4v
wG82UcCk1+b+0UCXKk6fILPaSZd34ak4P0t7d00O/RDMMwTiq0NarmWJz68cr3C5PTGbOYSFIsJJ
LWilG0/79dbo8mffrB/QrKnZKnvcBsRyoLoonHK0y7GP4a55gEAz9UV2oBYMs/CSt9VJFVq4TS82
A2vy6cBKtspRJotAjAZ2zcPwGl7uzUpJOLviN6GRhdhx0htv+xnkJWTxh0/gT8/B3dFqC7Z327Yr
HeXfI7ype68eXbUtAix4lF6eVaQCtbh67BQyYB0BFIbBQ8mHYexh//ZbBRM4ZYB1XjAYKqhZRALN
N9WXHwhYSRuk6739p8vsv5nquUxA/hR93g4xz0hvDjXXSENDvQCZSS5aB7AadTYPdElTHTmMQOZ8
2lw4+LTqofDyTghj61Fmen4rgzV8/xp25NnBiiXVno5QENG9ZT6GNhvRK3OnrWyu7sYe9epwYrQn
f1uyoApFYiL+Y4k+WHxqebUccmR8GfOHCr9QhMxu3BCc0uN2NOkYzdjht5LNHXUELhqf+RUlHIcm
Q6PTEzgGwhZOoLXoXwneaL8d0t5B2q8kHpMOVStQ6Fr8lP9SfwFTICVRhFzgBoyTCORAAXPlBY8+
+Iw60NsSIhmUE21+titoCBzbbCswIo6ButIf2Q/gjkXlZ/2HLjBhuMJuDl7eBsoViyCU2MHpsqeS
wRCv9hxcy7Pj8benKw5th0FnFZjxPEjnBY4uyfDoaHhbXt41uBXRaXDY0OyWZPZq/Y3bPqB8Px8e
yslDswW0rfJShL0DJHTw1gSXuc2Zk4V7SnMPgqyuof2Wezj89WyT1Hmb83FdkKnto2GQtVcGBxvb
WBL6kSuVwliGNZthgEWv1zc+YagDUoY02Fq5lp4rjVHt6N2xRj1+2zImPwWIDgobcAADFt5HCLFp
Bp51vmRLt5BX4tlnxVSHbBPo0wJBs+3ASlzU90RazuJhUoS19qfNfgBQ4tutr9kBtLqJ+4YuBR8l
WGAy5z4hF9WDSKg8KMwK4pVxGvLjoBYmGRvh+eK8eNp1rzYhYcGWi/I97kUdLBescA1KBgqQt8nB
Q9KWWXxo6Cw+Izvs1Pe8JxOt9pwE1+Kk5SPt0cbyY17vqxQ9HLErgNPgw5yGqPDMaVmYxxmPkAqg
p5nE52Zv+2bVDXnsA8SCMV6Yp9PxistD/dye41r7VEsPsJa771YdbrkbelZPYl0psRCQcPKOn3NI
yprrCqlqYxmjbmuavEQ0l6dUlIMJE1t3Rr9t2xh9L+d5ZbyyZ1oX0PQSQG3R2gNL1om3TRXku40w
7PdUuZOfLhAwacTZOW10cslAPa9Ppiy2cXBgqUxqnrYgKWr4HBE5FU8NDpbStPeomrEshNZ1OmHz
4Joz2EcOzdWe0hb9zIRgdPCKPEqpS7ZyPJMyL2ZnpQNRqKvDbxy4IW8rCVs7xvB2VXp1z9eXR5qW
o4Tch3YcRSXUlLijgu7/mAKhrsy4sva3uf8usUID9+o2KZekLlMNf542aDtdVkYAKJvxUB6i+HqR
6JMLtLk47PNH9z62xAw3FdMS1aq5kirAs+5AYFGh3SC9IPkgYUA6XipoefXJhkHO9DS3o4khtBNN
C2Eg8CKBfNKMpT/wpo2QfIAW5mhmm6NlwoC5KTYIOFcvIXRNLxkE2e8AxhrMsjmBT3bXbDPAhmSP
+7+CqmdmZ8j5vWh/kZHwSDl1IY6/xZYpbTxnC0FnS0soShpa6X0cs8KOB6gu+egtOx7VPjF4bcjk
uTQWp/eY5nxQkLlXz9JAqzwwQHA0ytPRgh1cVs0Gootfw/lMnxoe8gDkaoLajDKsVlFSkHOBP1ty
yFS2Bt0ZTH8VQ/AmWgeZ3/8tfmXZcUYDVnrPDETNGjWaBFrUA+MMEGl+IKaTWoViSWmd01CAtTh4
v7Z//wYGcurRj48EXlZHkJpPpyQO1T+ThpXSvDzsLRTDDyMLJ4lFYjcNgAPCZi5qzVoXgLNZFfwe
Pg5TypXHXRNt5QcQsl4D84siECeLKL3jIvJ6i6aZt/Bny0H1TcO+eVWC9QVqXu2UF+nRQVlFGV1r
EHg9Lxi7rO7yMpF2306BoDzAMDXTt7s0TyR+KdwZ4BMnOXsgiKKxPvw0YzhN0wxr24v0ilX+/2Wv
oDiPhwMCq4YyNAMIXKrruXm6+43aMPfzbQRpUfyqaKNtEOj0lIbGYltun202JMksVyY7AvZsNjTR
u1k9Lxibd3Hk4xsMl4oVmuh7nr3dTbA8t1ZDpPhe6OhI8SNq15szBESzNG5faxQFZS+H24ZxvSIJ
xdY+YjJlVl1Z4cqRgfSorX7lO6DN0KD+SbWoQ84gktBSwfkJfDeWXjcoElCx6RzrTtgkVYaA7mAm
8xkUkvmUWuGVA0BIbdUrRHQ1e1RMNneRlijPtue8YedhGdZn2wjreSqQEh8m/OjP+ExKNfLn1/6q
zpTgT+vUM73r0hhMjtQHT2t3O/fDuIWmVHgo/ljPd+MmI4cvlY+LHQLd1Z3aCKEsR0s/jVRy/c1g
yoOwyfISCl0R6pa3Ot1gHqx1/CYYoM63+ukUmfdeQCvvcpRfsMCVmEHa0JUT2M9mr4aM1Rpbx+UM
Kc87OB7mau2nkpa4sxn4soT6UgYgrXFeg7V6Hd7IFv1lg0kJl8cRLmzv9XHa6tFfUNQiZ5KrlA66
GJSF/Kh+jYBfF2/ySJtOOhPkD8wmCtt60wkhRlKN+pk6YXcxmtRt7IgMTG16Fy8PdrgOCKzoJntN
8U4JbwBbZ1zb8C7r6FCYavUVfeG7auMoPCOyLplLYtxSjP1j/4CbbtQhpOum6BnKRiloPVbpcKx5
n3Y2GCqaqGJzeIlEdkA4dbO7DQIityMsYkxqEsc+wqlC/w9zJPcWqZtEw7KQZDFYOx3TVAFnP4jV
80Vo4ZeSxVN/LKEA626dYE9mKlRvt+j220zGoJ0RrS7yCs2dd/dt3F0t1YMVlkYPTZy9yopHTdAU
FRCzhvKRBgKwV0gCD7WMmxvq6oM14nggsLPzr1QlBbKn34Drn8a3c5KmwTC0LQZ2qQH0StJvwgZL
Vdss0P0LtT0BaTYpRcIWOTngvJcq+yjkpgWW0Wuxm4c2R5WIk0m9fOI6NCjmDTfs4QmaVEUmAD5w
jbOhExz4oBHHC5PWHqWVGHv4xNeZutHoiMzBaRj4AHtYxbzSE134scZzIOMqdfFxZx2fBukpuFS5
3e9vX5STh2/M+Au/8yrCGGihyJH/iNKaCdazwoMQhlmJ1VvclV9lwsPbQbn0JWvq0s9MTNCG2pJa
JnXmP5GaFc2Lc8HdD2q66+mQ0D9Cte46mKWrXMpYU8W8/NlZkLM/HxoGY+fDVqQ34X8xpze3i0XZ
e8+M/j6ADsnyRrLt7j/uvOCV7g82QWHaY5xkWevuW/KOHywbLc2pZq2sjJQ96HeiRygF7URRqtnQ
id2ElE7kjT/zT6OPg/Hj3TtgqDuMVMs6wW+UI0fAZcSuG7o7FuHRQ0JliML8MnYgz0o7W1CkFQZo
xsxSmRiFEwKg+psgEHlkHC/9UylFcH24QQj4Eiy73bWFKSTabjCetLZjh4uCzwGtY1ZexwxipldP
o5ZwgXuk7r/z1gCviSUMW2z1lX6V+Yz5UjI6GDbNtqSVLiXw9OohN2VtxI8ff0fKtT+QtPufEMpA
BkgVAb9UlRFuACs3j/JrDb5Kkf5a+TAHgJv4mncAdiXHPBsBWBaXszMFauEuBKyM2C70E7wYEKa5
ricHwNAyHNeWYecpJjvX4QLDtA8gZH848LnRfOxHoVzxpX42R5ZHGl5unFaqKzOdISOl5faomYGA
0aiQ0+4a/hgFPAJalPh4LyG4p79FZK/HCEUY3XeMvjKEuV4X1h9lXANo3OyIrD7m0rP6B2kVM/hv
aB/n2Fz491vczuDztSOj3Yixg2rhZs40m1y94P1nbh2UNwLJhS0N2Xv3CIBByrwlpFZqAE+uDl5K
eYoOpkV5KyY3LLxejQXR1yOkMmFbqaEVaqePyuqvLfpYJelhaLYJSIV+SmfD9BQaFpW0gbVNxGS4
rUwE6b3btgaU7zIp0FTLAmuo77sAVNfGCOyRX7UJCsOLKsWLAWgyq1V2w+ce1EpG42hQqTRIXVhU
xZkrtzLx91opTxdwNPAlzQDavHwI/guiECp24IWsJrrPKRt8F6kAwa+pWUExqp/7BTpqs820DMCk
AvgOR3OQKe7k86W6BMP1s+ea7+fx6fHiYq4YBQv8tLIE7niPZXLhGSi+q/8USLNp4DsItu3Jdzlo
wTgZHxMOkUGMz/fG8CiYaghsGHVWDqL7C5yaZAr9Rxv6somKzaJ3oFYvuKrFpRT2xDlSkI9Weasq
njtJlVJNNiQViwN4tlG/tJvsVbrT4dPKtSHbKIXu2rYOMhxvlamgDkn20G0Lxvg5bQcgnQYi9jdf
4BJYHAB9aXGITFX5jeH/z7RjrXwYGgkBOZGF+YUB+4H7ViEszgWqe5H+7jJVSovoIc248RnwZbJV
DrieYnQG+kfSzY+N8T1gvvp2iR9CQpyX9gKGTaLzA/2kkTsRcPPTYB4MBpL/ifYQQLgKp6wg4Lo6
UNP6J7zdtou054JWuBh7JrKGWMllMg843cra1U7QeYUsbb/NVqxxzOwEnf0XbJXOukeAm/jJ4zhc
SJ4Bo3xfbOLUJHPP4eGMACmIAeI5kxqsTzbOFA1MROoP/by6owfB2txtgvKlB/zCO4pT47vXm/qp
MQKd6Ek5CqQcpBJHegZ3kbiTbeplhYKLJEeRY7FXn0IO16eLD8+/IT7oxkaRTxq3/8xdmmT2L5xr
rvgAqoim3ZM2awHQkLkKRSUIvLTAeO2zL74/qkOUrGKiwt2J8qz3SvkQYmrRXU56hyC+EDVGnDWq
Xfgqd//CHH99eE8J5msvA7AvOYYvcZX36ME3y0Yv3SJcc3DOdTUSPTlZ390f44Os8XHzq/HNTGJl
mkfVmVsKs8UH+3Bsp8SCTcL8zSXAl3D2JJV5HlOKpcrJwlbHZDElMt+deRasXm9X0C5XGXARgPB2
ePxJEIi52ZV0EAYEhpf767eE1j+OuCxz/fD/ef0fjWAnvfWGaZGwLT18Vw/x7QViDGPty2NyNirr
Cz1VHXsj9AO9S9LisQvSy3PyOHphiBAcwgfJ+hdcWq/C3rQLWK9DBLNUwnPGYjmM56B+kp6etEbP
0XrRLE8WrcHBxxD6eObBJxurg1Q+c8v36r+4mCwU+UIitkeurUm4dbAhiCSsagZ6xm0TuJ16EnWO
wDfe9FsXD/0qdRnPzcsW+FUi3CRjVZd8y/85Osnw9pNiPAOZYUV2JsQE7tB3ygyR0n2DT+w/eSWO
GmS6IuXLJoo16KM5wtN36drger21fxkdxvjQz2QbNkhX45jMQ944RzAbjZ+hId4BtGTbp3nWzwf4
DtW2cOCghbTbPIdtk+VmtzvcLJKFphin9/CO0Ps1Zn8ReAw1GGAD4nJ8TTwiWUUcWfYGDVHKz2A/
/Wv4KcuEPJ6TwvsxdH1JP3Nnv1P11E38EOZBa1skMisVyPQXtoBoIKuguiC+AYgr4KPA7pPJzqfP
7xVqqCDQFnhr1TLAuuC3yR73YUdGdqn/YQ1mjDgKmUi+MwAsftUVGU3VP5MJL5EcxRsEQnh3Mgy6
pv0zBzh1blht7JSIVgosCFkkdaYiyMgutfcL4/etv5vOBnQ7ULDK/S/FyYkWp6JG7QlcuV0PgEMF
6XCVaCJdOXVS+gmBHOYH39PFnTSSxCwNSMEYp5m3P0HmdpuJEEDubsw6ofTooAL3/ftIolIRjFnX
+Ps5ObmIRmoOyKXnq201IQKXuATbL8HoAeomKrPNRBa2OKfzG91Wx2tEjXTshxi9zy+Ra49oIVQq
DVEhbj2RpYJKt1xZ8EAErO+ApIDMBcfXhNBHr0bifwTnI05ghzmkzpzfnR+CpxkN+yht8lFlufti
rI+0uKLimYMM8KD6K9OZE3iolvSoJBBG72ER+a/fcYJqz2/enoQRIKAL/j+nMIXqgy7p/ic9dOSG
zQ796Hv7Sj6VotE7Nsh/DqgZI1JqGPc6+0jEcAb6atNzafEc3Y4XZXrIibUlLpbSxDbSU+GybBAR
zuCxK3xG0kf3L2tjsDENddrr18Ck2rd2W8dLdIfvurQGzFU3dqdTEZAFNptG8eQ+/f0ze9/VTQjm
Xtukp7Sr43KNv39SWGI9jjItB6Dq/J4PGiDbE2XuPdkM1omBN+BHaQ/u1corn/M+P5GLqd80rkHC
C4OiYSYy4yTtjlBg8l/0NxfIMeropSLZ9i22ipNrxounKXiFvechPa017fN6Uz1AiULTekPvUauc
8rL9Kf0ruXoSEyUG6xTSVTzCH0ZwOtCFFIP06uzc3kqj64ozS7W7w0U1R5+/5wdGkarlMqeU8QQ3
cCAzmW4ay/h24UZzJFd4jgFDuAaQQvI8jhJrJaKwJUsxJvTjYAUJ2kcdv4BvX5ckIPdrsG7/17t0
e/OqOoDAEFOtW7ov43VkLDFyatv9oX9sWYfQIhoV6Sv9WAq7eRzopPy0KvR86AtAXQA+RP4kOvUg
Ouai8728HSDjRWHIdveiYJHoO2V3WY0vPxaEV+VbHjzLlbb5KT45Z7abGBe7T1/NxReme1b/9xKn
27J4ve697LPzduPdLFW2tM9qUfjg4pAXQKJvqpQnpVTIMG9WGLA0SUO91EncXvdFARA3ZU0v30b+
pi78xbcgORTNITf+28G5zFZVd8hRb+YsJgKX3HefP5x4mkOxIy91a8HUwgd00D8sN6IhSAfViCUm
xnd27aiau2kGHtO9V2mY0cFWp8r/GqlXcKPS+sK6SLc2zovWzXBvMthvFCzMoRywymB6pzTUvOxj
PaT76iZRCfdiDu9Dv0hF3cdTmeX59bfBULTfIFWc9gpSfqF5TGR4vBn3/7QOlNreMVfQUTzeIXZ7
POFB5NbevExtKSqrQEig2gSskycFr/F+0jVuZCdORWExrsw1aSFe+oNJShIVTpyjG7I5g9t+P+aR
3rRxemQKHghawVz8cRjG/+hCfdQf3QxW1nFUWZ4JP6A4j1IhmE3Imv0G60LjdGkLD6zT2TqeX/O/
lgQg0TfVnVFXnUR5j4uOrUrn/IXb44Qi+cudM5FV0tCxRBNke8YnqHv8IghvHezy5m1tAepDdlGg
9hlwVEl/dcwwOpVorUjQEOzMc30kl4tFH52+miD/JrVn67Dw62P0r/18I8sid+WCEzwUJW/eJhgV
Z82RTjaAlb5Ljj5prOQK47up+qqQ5LQZ83DwZzja5jDMi31E9mtVAgPOsz7llcJ4TqV8eY505YPf
oarkU+cT13sEkxBZyEXDOcoPgdEuLLbmkskpdPjvRyBAvB3HRtAxQqM/GoKHLjxwE5YBGhN+3ShA
aZQhvhHpKfZFUanarGOVFzYI27ieniM83+/EVfo8Cl8r3P4QEGFKFf67TT4290DXaVuqu6XwejAy
pVX8Zfx/OwrDR9ynoca3iUU8Z9kv8EEmxlaMUfQ5/4qZN/rD+g9lGV5Chxn+eyzzucXrY57ipYct
/T5sbfI4uphGzKlHywNM75lXwAOJxZgWq1yzbKQvPdYbbhZ6h2ArujON8ggYn2p5qcmHzaNv5Ef5
nKx0cXN1PwBSIMvpLUW5YNMY4guYqCRrl+5+gdoiCOtGRbv5jrXFsEXug3OHMwATBcYdP4JuUw2N
1uhzlF43Myhk6HxrJ9I1FLoBkgphKUFfLSxp1O2SySjOv/ssD93U3GW7QiJNH9Ym0ThLYJsPNVNy
/rtMoBESVl+urMZOmKL2zpjGa4CuiId1IJwcaASU2e6tw57eoTekjiBpsP69rdFbUTW6yCzyCp4H
5wapn4mADz+E8fXG3QR9xNlm6m5pNgwzNS+cYtGp0CHVrbHcWYCY+vuWNtOrdCmHzNI66Lbjwbsa
V53mJht738UbsxL4oXypM6WMo4PQvTA0+SxYeJvHQaZkozd6Qfu5mHfJTMP7Ogsb5713gwDe+j8e
cPG7pAJ21uLCFyro92RzbDl1uJRu1vnXVUHBT/ek6U4vI0Se6r7VLnOfLdYF3pG8LEtj9XgTRmkA
CChTFvJCyq13I52MXzrCKaycTGcaUtoAeZy1cZDsA9T7DuW+FXYJ2p+68tHu/XiKIE85lMiYOuCN
w1jIw0ohZ0uTB9KrN2JaFycJznw3kcE5vCW9xKGoa0fCFSH3DaOyMR6EBDOTwhLEfzk7EAUGp6Xe
LE7A7AXQ7z2IzXDYcLmkotB2ylbpvSzxSdtCL4dw6a4/H4frduyAXWsVA/4SPmy54U9vnJf4zb1G
nLMp+47FDpHAMmdzx7Xt9p99PUNTk5QzElgcUOJhDucRf3ROMJLrkklYOfCoX5WX0Dbi1KYF8cFL
zb700WdgTG4k0Vbdd8a2NL/mA2wq2iZzQb1TdQ3+ggZB51/9PB74gDmX3ZZosZEvA5xOfPGJtWI3
j9l+73hXdPh8lq6sg6z+kuTKoQzPN6c7yZCTN53UhigjEcxu4ykKzhTN0aIMyt7vs/t3EwAHC6av
Hc2xJpg75/hvXljumplwHa4H0DZqbxkEvkBz7h/T4i8IXW3KNt/88LA5sIU9+PQshNqfCESMJVoc
irv9eC4nzNg3qIJB33lzMsg7I+h2AKLJxgAnn1ek6fZTkqvG5W0iFYZ2J3naWiy0DK0tviYyQypd
AeZY5XRegUNZuUhXbYSYpgDTLLKruQ+JjrENJgnND0x1S3MnRfybWc0jlswvnF/Hq+PeQw4vlsjD
PLYYA9TkcggzjN9xO7xWbGpEx1mjM3opU+OphaRY215mT50eLiWHVFcWOxbgwqFOVdY6jegN/cnH
MSRiyr/1gMcx6U6N3ROcIKahteL7eGS8bVzBXD7Tl7PAMUPX+R5kOdGAWwsmbDubq6Gqci9LjqJw
4m/+JGUdoFl9QQDPlaKT7g1mbQha7ClbCebKTldxsxWVhKWxG3tFQl1qFMg+pUnmvLcIGIc1c8+U
WOmFI5DasbsURpf43LZ9r/gtqh+Vt+jV0zBthZbwEYU+kN6Z9ZOUApIMMpAQwNzwP3fbmNbJ3wi0
o2bnabhRizTMHQogDtdm4jQLDpsuTxuAG3NBTugYCiS4owOI5133ITCkL6e0vlnnvJqu84/BpspD
XYFpsFZ4ZTh5rocTXWpv76qF9KA1sYTx4qw/+E0Y2st0+qb4vRt+9ZgEOP1uxRB0FWrgPOFBs01r
45OZQhS4HQIHbEXlgz3CZAE2HColUNx0vrp22ky5wR0JtJJJtJ6C4jRW0squfuCL8VPiyhLdg6YA
3u0X4EXloMJ50luVIw/xO4dgFiQHwlUTdS5/ySDJy9OHeaUUTl9yzLeORgeaFS0kvq0C9ynQI8tc
ACORm+mS+VbbjKgQ091DXefUEgex0lRZ91UcvByT+bRJoiWQBTCA1C+8TRuykyKAsFna+nHgj1Tl
nTLmH3g3YAnhTdkZcVMVumXRVcpcFPQB30KRpWxQ3y4zNXIgbn+LFSh69PJ7dNqioaYKdj9/xD+H
p2oqRa4fJBbkG43+Ouo0Kaoi9mdGJhVszARK0tuMJo+jHh2GSlqWNxB+A9DOo1gL6+O3Mt+feFPB
BJPhfisH9MDMPqCLeLZ4bF3aytPad4X7t9g/EyD+CVS3+bZkIjF2AJSErdanlkAWvyqNFlwJw6VW
0ozhi25jf39UtD8nHc2SEtp+/3T/Nq8yLgemz/um3kzK/UZfON6pKiJhjmhmjP1wlfUnnUyld92k
cy3zfS2vc4anheMiFJokAlmMvEDKL0m4oO4GjP6dy/CQBm92zLDjkuLv/TBfIt1BJWeIvAqclqr4
bmIRde28My54dXcHsuWGQoqtGhBtB27VCJIXGqBf1ZPdeo3sKwd085RrD58YllU8dvxgQU4vUfWs
MiV6CbHrIfRP7fWA+j1PAtTntuBgI23CY+jhyCu1Ch2WdCfOQyxFdZ3K2TR4aHTAgOVYrIWMM/vK
AFWMPTi4jys5dGBj2U4A2Bhy/9uKqAJmyol7Ez30cyjfoDAIhgnnLlFhfljJRQaclP+Csz3AQX8/
rzefu36esVXctZXb7WdcMJxIkaE96PdPrljfrvXad3+O7LlV/5iBoJ3M+1zfdAKaOSi75pm245Bz
icBHnIasqANZ5CyiQJDm575QabQIyA9cs0sct2Nqbzky8ObolOjhXgpnk58yUiW89o71y1Ero9SO
kUkCfZCXk0X7aPTv4MW1I5IUv0rud5IcpITFG0yXamBm0ozjfwmPTD/bMunf0LB5e7lxNuaMqfYg
YjobEWuYYCfyS5zXOaza+l0Dp2/nc7O+6j4BLfzpYSmCDzaHXEFzOgpD2Ro4B/iimtL3yUWs6ctx
bB+LrYyh2RT3VrCgFX3U+/dLxCJP92Cbnvz83FPeJlAL8/5ZpuiWbZ/mX+Haog4JSiBRx3o+oLIe
nuGpVyHpjo4XVxyVHx0FqoOKs90lrlfl5zYWX+ec/zAVu50uU54V86ipnkyJyiA/mrnI8WMql1S9
aSc6Wl5mUGZl7fUrt6VV665avO1DS15LCLrNilV2gr87akv5AgVw+Ge5Odd7nPn3SiYpIe1JnKGe
KyhcqIVsEU+WI66l8lyw8F1dtTZr22wv49sbysX/QeShpondGGlFN5WXClfmbpX3S8gDnZSb4pvm
U1dPp2RKeEdotdgx35D+xFO0KtazoJgC6IoqB+74f8bsPe02NtB5qwuzw93RTwBfNg1vK76mQ95O
7gLjYesIf2SXsYGzeDPtS+ZkMwsS4XBOxDekjspo9/brJhve4lGhKBxsCDST3RTs79a7TRSlK/Pr
6dRFnQi2tbJunircBnoY6yfQduoyewDRBoGqEktypKe6LBVrY50tWwD3K9l7YtSAgIjGSJJIlrRD
eRbjo+X36IlfcgcdQ0f4+UKsXnPKUOHSFiGr+hSi5yUlZcJPRsgGxwqnXiy68v8C4UxO3mfNKAdQ
eCFckkPs5nySS9ivNeBj1ZuvLY4YgJrI2mpdtaQEefX94UsPQwexEvoZq62m7MWbIufNouhiXqJO
fNS3IRtBfOrVKUiNzJcBYcCQkX6PSZJ2/IDGsCl8mbUGWsfM0lih51TNif4HjTTKC7uoK8fDfNSx
zDJFP4SHbAwTyaz4rSG2Or9MDbSRF+pq0U8GLtyvctSA1Aus/sLZa0G+2tyC2t3jI4mCJqSjS6dY
XEMHWtUU40VcA4SEeJUj1+coFma9JKx5MzvxUZMlrYng4c9d+73ZR05tgMycdWVKomDRIOBackqN
grBq12thyWyqpawEXgw1cnS40DYppssORmOpXDt4ix9QILyuwXYE0KjJ52zwlGdFqigNNGHqbPis
4JpMKaTcoNPMt6gy8POzOBWE/j7Wtfvem4dFXL9q7x/sn+OtXIMQ/73xSG3wAbp6EtJ8Eu48vxCY
MtvimCV2KptM+iQHdzieBLaSpzVIq8U6U04sdXitgmXYslUI/w4CSw524zFnIjri0A7tSZP2+QZq
+nVfToGoY7JvTPGDuhqIMk5UGkGTFUw8l8r2tjvujXxr9TE06yzlJXUMnNuoLXgsus/MqFuwRRlX
Dd+FjcjxQskNrAldV2MZGoGSDZwx0zJwQqtBZj/kz4QPPC6lqkDE12i0zIhUjTrX924y9odpmsCu
CPs79EEn6wQr7uQ+EKbGmbCn2HRo9JWPs0pV3nWBzDOXOauXOadjc6UyLjwTJOsl4J6N7x5zHTxF
ArDXAHOq8zHfuDkMfqBHn3azXdNb+mUYbpMoGZigfLNuTgrqvUok2YaIqf+zvu5wlePYAEhDgJRY
SyusudkE2qItMV/7lZxqY+H5mhC7p0+AhohASBxX5mY/T5FY07qI3H+38agALIEg2hGqc8K0Zb/l
pR9iSybVIcIFnSe33fEpraPGKkB4NWxaPBjcyhp5Cj7VeCrb1mdTTuTJaCIj875AxiyOL65mZ1tE
oxhhd43eES7mLJCC39rG0rxGMSMq3Ud3NqCb5u070vVr19zqmhsELv37m0ejlvr1CQITfIegBNcB
Bxo/zWGFZUBY3TRtdL8xqiFGzAxlCdLPnkqy5aHUKARpyZcfsJvUNr3lj3R/1ggYFe5sCMCOvjIi
MfwYR3lcu96b6A1kgx6fTGWVIVgRWhSaQXTqKC/28dkySsUHhycvxGRjbM7ipweXgpLQqpLdl/oI
kn+u56wI7TOsKVKMz2sviXJ6mHMHG1YJBku3Ujhdgh01LgSJK/GtrPdwDGJJ0uy5f64sbZEpkIPk
zyHCugF9m+Wsn5Yt3T8oRdmA5EsJ0r3mc4G6XOwWP+lEoFjz62yL3Y6WDJ2O13CrvSTVwewt3Cat
IW4UD0N6pn0skKLNqzPwNGBk9KVl84fGOnzvlhxAOlmRPugvXTIlgMOE7OICENv01Orr0RLSb7Hq
2/78k8kXIn6NFVEc/TPA4aTcemDGex2QDowUGiowwim7e1s42aRKI4PBoYLsn/0TZP+u/OFJ3rmU
3u52K3H9Yauvs29siA0Cqh3DUlgDGlBW9mvns0YunXDIjlFmwVk3ow+Hidcgsf4jkKSa44BvW8ZL
e3dXFH+OatebE+0T7iv16wLcMHEjg8Qj5VHoDTV10lt/81qtc0h5xgk/La/eSTJsKZG0Qz5tb8dO
YRi1gpQ8lk7aYAyzEYUX2JOvaSuNn9/il7wMY8Is0V5IGIcHTI0OyG46jwDmF+kIAp0Ai95jZanQ
hc/gkdaXGAh7tlD4c56UsS78dGLFGrCK+9gtReH3Lk2Kb2DvDNU/83mhjl5loC5idJt/0OgtdnW2
s1Z22uRlluZ+wNRGOi++s+r9dr/PEDV7KOl/1lY+0oEeE38kWC2i8CJub1SFAl+c/0sEutQr18l9
Eyh5235PMMtYn9T82DsPFadGCnA2qQR97TfRqySDA7Vk02te+f4LUguo1ytOXF1YMou9i6QejuMT
vzPIGS6RJqzAstYDHhr98FcrUZUwCwtNWZbXYiNDcbJ+UnkQQI8O2d0HMG+NEplnWioWvtAnPws6
gUeKWEkjRmndUrnnUaRKcpAj8JMrEbMQdDzFTRE+YBGkeMADkqw7aE1Ke4FMt2f9cKDUBazoPmhI
lOi7z5lioR5Czxbbqn51TovQhs6D3lP818vr1NkbOud3slM33D5+E/jAf83Bc/4CS5XncngINYCx
IDxrQh8SMoitOBvDcl3qYViImMt6yxCXjoHF7vqXJn2YA2z9LJy7W39HYGWq8WDCP8hccJ1NqvcX
Cq78GU+VQOoNRBY+CKrrIFeZ+5jTA3Ntu/QMve7xV1NvZKPC1fOaGPZN0SKz+I3OIi3L0Ib5ttWy
wR8XRT/jDr0HRLNFGU4J4giUSnKuy2oJtMzcB9+qVb4G5sGp/Z3FjD9mOU/PR0ido95bzdFqbzPP
ZBWgZs2G/xix1YYcqkid1KdGoucc+9UwU7UClEDm/3RnQ85Jf7Ld9+uadb4NE6hm/cTmxuBt483F
ZTmkFC20LiPSXeNT6oShihegl86OJV/9NCofhtJPAls2pFHE1gdlo4kmh3YUYxkR5thmu07CfF03
qDooVX1L4bwbcdrmpiDk+5O454ertaUSs27tDmgF5B+U4sIAerc/2mt0mI8DWZ36sCzRtJa8Ucvz
PfPPMrbcimC8Ove69T8ZG8lSBukkAq/mOo1ODQe9orIuEcasHTbway6HPdbPVDZf1kcLzpNfcBiS
7Kp4O/io74OKT7Z0WLmx6vTJk+EiBPmol71OJ2TtrVtguBzF/XqwH+8yPJuabpqUQApXXqridv5M
iERUpyJitQyKVhWfLutUXbgzEXBibubEoGpU+jrIjUCfpaFfKvJfsqGHpfe5LF/Izb3GCnTv26dT
Thaf9XOLo7Wep6RACC7J5ETRmdvThzzhVOKmiVv5/F6QQJ3Hwluxwk91dqEy8AO+x6LNktTxLpKJ
QOLfdvxMSsYwtEQ18E+lnYxlljFFoKwXHbZ6fEuxHb1bfUYT+ag3hVTFm2AZVwVjiWMGsV8D2vAZ
CsVuf7CixFC0WiVI5k5rd7+RG7kX5CecUp+IKoCxKV58oxL07b12Vd0NnTufldby3ui8L/mucmZe
WkAo4gdB9nJ2OiOoVoIwASfuOD4wFjxeB8b/sBlF6Sf6fa+6r02GxuooTEU5v/3y8GInst6leCf/
O3FnK2AWu6kNPq/hUvkRmA9qhrogxNlwjA5TfraE3HAQjjTNib6MdSKf8cofpX14COPUBMQddvmp
QMJh1WeHRDz9ramUW6BUBIJVZb5kAxvwPOt5kCmNPBV73FgslBNYW835DrftZnBg7VgRI9Hy4Ay2
Ac85cycx8WmVRSsGxCzDu0MgDktDAIJMXMYIGxX+c4g0XGHQqD+Yn4iB+FXXJ16WD5hy7cU7PF/U
oeKVDzHR41uHvOLbMgGsSGd72XWO5G4sj2xCFja0Ok0ZVpMPPmARjt7vnTFGnZz6hydC1nYxnB7A
SQ/2E4XuWuIP/hKKlnHrsxfdM9m+7+W5YfYr85lsF835Jru50zI5z1RH4Ss7Vnit0kWnQZlWkDVN
gDnjY1fcnDIJYwRkHoA9CsQHGjT4CVxzZBgfuQMblmGGCTpvBnXRxOPLoUhTfUGKPEbKfYuepI/g
WzCeEcjqLvkNwfAqTNxZWgzNYmdCyLp/qHsRgYZLB8z57lNDu/oY363T2Rn9uvg0AfFAHfQ53iH/
QGVa8+lsc1Y8yorvIBYFZM/lL38J585aztXkZtrYXqsRGjv/YhjcBoIHmL+RPduHqOt3BjwP8AYi
yQ1upmzGs3dLysddfe4nzVTDJxBADMpEe7X+hCzUg39+Moy1XvV/8kRNprPkYFq5V4S82YYjXlIG
1RzhwweS+2uQWQyCb+PXTS0YKTxVzGMx5EleGr1HgnkTbY2i1iHODucaN9N0I5XVZ8HxPcubYD56
kKxiPqo0/RpdKfQ1Zp8quT3z1aO9boe5ggZlPgiTs/KT+dFFZAEqueNscNio8a1RLpvxQ4F5WHIh
XnXUZJ227+QFj3qFccM2jSL8n+JJr9Z1ObNDKtBJPTRwYK+Yr1HnCpVtBZZO3kv8t9yhuAaZBqeM
C55N91jWio8RqWGZLJGCmvmqyt9xBehFRcDkZEaBAREdrNCSPGydn4m5Jxy0LbL770q32OZqC4jW
fSLa0IQVrNx0jIVjiED9JwGNq+YhE6szMfxtvPKtd5CkwrwFzQRiSwZpOSWVZylPEuMwBuVUPFaI
JASuQSXwq1bx8TPaTirvcJxix757YpkrTo5qXxTsNVc9wI/7L6xr8yU6P9MvYkYsV7ZJDratwH7a
yASoxKAInZ8kCFD+3m1YNbOnsT0uY/EFk06Yhe206l9+sfio+L8K+JQF1JM8WZXBl5xnNAqeCHJy
Oa2KPQJIpLKOx+0HJHzTT1rmugPfmJM/OYybzkiKoddX2WuF/dfJby27wAy8rRYdjdl0rmXPxP6N
tXuzYxeLVcQy6k0Oi8Ir2vWOTzazkCyK8kXu3cg5Pi6TKP9DdQmX27PGTL5Ni0I0NYmW5gGesP/H
0nv2jQ2lOQyiu0NXvNcW+14lEKYYNsWk3Bsg+y3ew35nUwjVODTMBOryZD2x0ULqiOue1dr4zF0z
UbU5p+q+CgsfG4Ch/q+lWu1zS0kNgPG6cnf/igG/eNe0PJ9Qlx0FHxamTYyS8W01yYX8fTfspbnt
8pJgI4zrhKfPs6YEyLCa7dYnq1NAqvfhk7rhuZtoe7l2Qtk9j+9ooTjQdXNY9ZhACVTvC3zWp9/Q
tEECCvttR0icFWTGiTvzKKgw30NQROXUNyBlP/UgTBk9BG7Jt/3Pprgsq0KGQad2jyBcnqiKzSgR
uwq3dRjfrYiMXZPT3h2yekJ1rdsyMWrfd2hnsKRHraNBkdClsUoz282jaMKFbHNTNUQKHLwbkAhV
C32yqZ8hwCFjLiPuXRVTmERijEXsCZUHBTk/8XcJGNvjBM6ORNtJI3gzM6hkgdrfa7qKb1pHr8cX
BAV4ZWW4I4X4Jx3gPRUzqJacmzcdOZG2fWFSve+AyRzugif5Ud4GsvActKiNgB14CcdEOQm95n6X
UGEgqG1KiBmlhYOI82UiqgjEyMHE/4svjt7wonL6RHBT2p8wq9gCi0lX1l1yTtx9rPFTuRh814Nv
3/HRDUXy9+x+N1Jw4Kl4KLZknfxG+5QktNCJEbza4U5mEZwYFTPYk0N1B050I9H3ZgK2ZJ1ijC6i
bTy1Z+yKgngvUXV8o02A07iQhvHSoTZ03d3/sGKm4LxJSXuRTVY5O1t/SXxHMExDfUJxBoxzQyEH
tpVGXe3VTL4t5TdYHR7d8Du0npRBkD9ityiBdkq8LCyMJOAztd9IjEeGvFcHa3QFY8jHCErARTNP
dnLMnQ2ALnIOmHzeUz5Pnvlg9vGY6EIO7D9BmIVQRFmJ68ZDT+75gnYayYSETD7BMWpItkgn4Gyj
U8ojH8hWn0fLrtn2JNyrByBFBB7jlM9yg/ggCY2D+7IxZIVFC/31ynB28xv9qylVEk/dfpD04d71
3rG8HFTirQs275lKKOe0MVB6LEG9wBe73hh6NwJdLYryt0r0jc2l4Nl2SFyILMDbNDY7DBEgK4OU
6yRQSvlGfWq0Utwa9h97wQJIa4GnBSMn+4vdf3VKmKg4l0fCy7YbQT8I7KEx/yBtY+fYyoe0zJYj
d5n31k2eJGhIyQTRtyPbLaH+bz1hgHBqp4ewHGoq+/DIG0hP0h+BiA8kIJz0wENcInY7vInZADKB
MBAdUQyYmP272wBiesbKi7Ryikm9GSKrrA8jMDpDanRKVSMfcGArLQHxyuhxaeh1kOkxAKfc1o1W
8BhLQvhR7VONo4pOXEchUjvxnxCYl48uvG/F/Osl+nx+pP8w9yas2OViHpYraWo8TFDg0mkaA8jS
sw/0KFGG3hsk01cSmMRYIOXmDV0inG8OmZo+p3/1uZW1LC7x49HAikh5kYK1B9tv9drsmfTKTi70
3ni72XPbI6GGihEvI99lWpcnvSoV7km8nPuPKxtSi/LzsPxdBnnfEVYOIEQdUy2svkJrof5PuvS+
UrOYBC4D5cVag9yvZhWc5oU4POfeX6ug5F0nOSdBbtxclhnb6KYvZpCGfJK58PAPrCwRjHGFlQ59
GERqC8fy1k+7AR2W6q3SUTVyPxORlPsXBf0mSn5dTpiXPiwGTkRXQ4cpvup6fVs2tG1brMRa15Oe
KMjtoe8vWu8Y+iBWgpP1jvUSmJhb+RGGeVlImnUVT6lcWfNsV8s5dQZjL91gVFsXNBX5XQMgxMMd
/JpWxsBYy3BENrgxrI+mvAwGg1XPBxfGUrtyXbMzPvADcm2I/h5CK46MIXU7dPMKWS1LwPjMxIP5
TyPv5td6Weyic+4ijUVs2xkFaAmHfsck6/GAYVTpU7wv+RV+zLyi5lSGkAuO4GzFGP+xQju/JD7t
nfgbZtF8TSWW4GkvmLzuKUimgC3YYUvxH+1MBOKrjAkhzKonwYPGaO9oG8kfufuHr+zG7Lm5Oe5s
o88tkDXKo+CM0xvrRzmooS6G4XDaxJuVRRL66d77FiOcMc9aht9IWgkgq9BFcNbMXMM1JGYmhESv
j937HhjL+15kAGE77kJSxP4VOjAza17pRN8lcNk5bVo5a92hw9qoH3IFiN1XMTy7lB1+f55S6qSJ
pO0+LOl5PcIVutPfngL+geWFTFJLcz20EJxNWlJ9AssOZwmu29r4eLwQwzpfUJALR6M07QjCFmjZ
3gwAeqNTJx29srWlWKwx5SRSbCSxDfFyRCYa6V734qAlXVSOXQ11T2pBAilDd1PrdDJ9fEDQxSYj
v55WPWfx07zYw+Y4qDQqUPTIdMdu8skrcoUsPCAA+p6yFJA0T7hiC72qEtKwMiOKOQ4WAFigWUHA
gcXgKY10OawB2KfdZyd5waACo5N6KEqoAgqf48UIQA739eESJSrdckIH69AdtXbcFSoJ3Wmc0fey
WogqDBh2a1nOjot4BK4GRXnZ6e8Tns+9kUvrpXkOaITi6PSUzwaK7m0tkq4oTRS8H9WN0hnj2CD0
jQqee50/VPRJYCQiGn6z5LoOBiJdUMnLW/rPGFSN/OIEPwZD+etfFqBnL/ebYXFXY4n4Vn/kg+l0
PKtOuRm+xwtqmKWiDEnmlb0JVYiOmqCdZJCh5IwI9xghlenD1q41JNajLrJMIqHBLpQ8KL6lJYz2
VZpRVAXpsRcDF9Skmo8J3XXUnrq17GEARYNv3L2Rgaeqnzd79mLTaqpmgPuozIiRRgcBJyVDgQI0
qsOhINlA+UmAputdwxLHXanNBEzY08SuKijlF+LXoqfEaTe+CNzrZ+odyu/gSOwkIiWn41YCbtr9
AYBkAHszf0oeAlzGEtSVc5zmBlJXPOA1ifoYRqbrmXVGESINAoqjUnSZn675N1TfPUUHTEa5B1V5
KmNJ3qCNkS9kZAGg+dTb4YMcvk9ybOapEM9jjUdWPkiok2+8HhBH8QaSj7nEX3Dm2Q8CYZEsPKxZ
V7EUwtEE2XXiSnX9FGy7WPxrzpTPOZkPTP1C5p8sPH33mANP6hAlENKNl1/ctCldJsC7plTXhTgO
sBA3c7qtGAyRIEagzhFWvWn5QNtpv9BBq4G6JmzajjJqDYttpwZNSJtNcKM3uzMppV8xICDwRzGs
h7iHtV9tRuiQFlgJRn9F+vdK0e8ySSyK/Co9AaVpmYsOldywHGCG6iWrepp5evvvn4PE859A19pC
wMEQbCbldDyytmSI7m35DcXW8JZd5hIwx2MOvL5y39R3D/svZv+xgdwa5RV2hkg16gcHromxbqEL
C94vj2qGhDFN3elQvC6eYgsEi8E/9JI23FXv0yBPlnWLwuE+Ag27SuIp5ZVzq4lssRrAKlA7tm1P
MQA6InzGki8hr4303QkzkWu00CXNByT6KrCEfcCAuUdEGB0pwiyevzHl3fFwMVlS6iQM21r3xfgu
1MTSxWr78skAzhZh3RAnAC1fUeWLo0OPHTfI9VapIXKUF4yE6ohmZ+bRV27+NCDqLKbtaTgHY9zk
O0akipev+9aDEdt9Gld7tAxYwniRx1DS1tjfc1C2x3TRofM0A6n7MPZntLSxm49Psq7BtkW6ShMh
F2gLxCjxU60ZKD272sTtGC1k5JCTxEtay0t22PNzb1NlU1oMCn0bS6uG2kxCL0DOkxQ+OeBMf/L8
x4kjhBfEeo72Y1Wb+ArQR3l9BylaCEh8WionTjXM4Avp/Wao5xUbXZaBlM2idz5t1ZPREBBfYc/1
z/C32iIhsfDSAo4OtYlXVKrsxJ4M5CAFMxWGjldhZRJTjz+BWcgBAflvSzuOmdiKce152jLUc69P
OEmc99sDomjvDv61yPXSBQ7jaLDWFmHCltgvCqGGuRI4SBeRWmWPuZKGVP4JWzsKuXG18VBOtDAb
SZR1s38K737nIf5X55I0225/eoIa4T/+tlpodMRpSew1yuN5mVqspq1VmR7+eEYRG1DqHO7TRnbr
X1uYfWHFoutzrjeOh73qD5jRKEGQfeAfRugf7bHwO2DscJkwYBQAei2zsnWeZCeHPrJi8P5ZYQPR
5SN7eZDWwn7gvSVLVHfNZEaNWjxbSYB8X4ixy9xje+d270wYjLoREEpUaVjJgcSjnCPSzBbxMIUn
dIazFSj10h49XkYRPxjEEdT2zVMG1FxYM9TiFBd2Jmf1ByJybVr3F63iRrmqQq84WdN7W1XdcJCu
UI3KzjUWbk+U58CGe2vMlLo7LfEquxm7PPH3jriCbustFGsOFIbJrHlX/0Bw2ThfAyU5aLzxJZkl
K/X5VRZ1ejDt/lGe7FZjDaEtF4LghXgSDD2DCNtAvESboDGX391091/jk1qIB3VkwsEW04U56MyW
U9wZH73Qc9ZsU0N/Ni7F9KsDExKeygJ5NGcJgDumHeWPRwb+jnjeV04mfcq9aRyW8arlvDNrZo0Y
3fRnlSk8Tyo3DDvyl9Etu/5vlbHajSHzb6awZNsDJW+qUa7YM2GSfNKPEGzTj0KqIjsp/RUYIBlH
rBlnl3z+CReSGszmItW4TKmdFF5Ws03szzveu50OzQbcBggBVsoLflN0TdDfm4wdU7KbmauR2ytA
zdaBF4Rlii7JLkKaXQHufVH6K8eYutQYIHtc3AwXVYuFzFBseb1DgJTTI/mu6HEhh7JdvDukjaD4
rp6e30upBDv3hw9Tygc7DJCjmjGxwFeJKrzHUo3JcWcUsVyiXz+LvF9fsAztkqnPcipjZ4DUpXRQ
SnYoBFqEybkgX/y8gUGexwmd76mwS2CHnyjL4YeMcVIX6kEwgr/v4e6+02d+xOXP0jJLyIrA+DsB
1zs7IsWETv6YyoJ9EdLyPjr6ugMe5vZR40qvwsXi1OJf2gRM/ADVNm9GhY+zcuXeZK5R1aDOHA+6
pQr8o36tJx5HFe4nmGZ2Ic6nb7lhUMPeT0koIVJCbQtmFOYEJDwULvtVTHf4pXV0bj2LF62AObf8
btSpobgebLQwSv9IT5uHcZ5+5D4exTQxp5teZnUsH/1jmWRPQru+MmHnBO0son2vknq6DeLQdSu1
saSP6CoOorBCvRy5ftWr1Qr2FnNzhqC5zXfoiy8X2xvIUo64HarFQImCHW6JMqwpMBpvLg3Wof6g
fnSGBRyIMUgSIjygxqlK0lQkGlnWRdD3ee/8f4Skm+Wb1Nt/r8REZnf5EjvT1kXdZQmohWTErMH5
Hq/9I8JyWaVJjY1R0VMMHjNO+UIGgsD1/d64lQSnFBb9cr6qVPfOqF22fGDDpvt5l7G6O+kItDyd
2TLuI4pxmVYt+EKka2OwNTrUSarU6ifMuek+e/bvFRJlMjMGH2FD1Ld+4wKlNyxuCGUrqRv8SJMX
lkvS+kBFVNF1C+xE59Cg08JtDoXeIY6kTDZvZuiWURkZZnI93X8sumhKsh9Ijox3xBD196Anqziz
+oNwKxD4kSt5SQvdorEHPWCzXj/Og3hh0/BG3O33bQtmk+stefhz+oNFXvyILGPkj8zbeaLGBY10
8WUoMcMHi0+xIzlCOnth+tGeSUONmlvwRLMjxP7b68zbRt8yYcqrEdqTbvtC2HzJQdd7hiO+zNPK
zbqtSsWxxqoA/2uZxYWOC2Y6gNzIQcyJA7w8P0JURJVpn7DKcXydUchT0sdrZBkfIQw2BEBlX3zT
nY2LzcBrcdvIGvUfMH2KnzXlZXw7dwHw5lF9Y+Qk1khmLF6BfPPBs+BQhfILxtjZ14TsuaUAkakp
UYExB4/6K/H9yko6jcTblZf6CKuXRUIx7IZ6hvqRIdGlCeO5ISYj3AunAzhBQ9Rp0k1y5BlOJPLZ
280Qx6wObLTEx/nxF/xKd3dv4T1zaZFwl5GC0tU8DU1QCbMAhEh8pfx8jFJnfNiwZmyJjhTlXozP
1WorxAuXe2xalNqJW1nfMsfiYw03GfgO115xZcgvLqNcLBbcMs547gEmfYsNlHqQWOwMv7ph7oen
yfW5+oNxO1mrfie5Xrq/IVlE8S9XDHPB/i+UFkKNUdpnaK8zKePyNrk0Oc/S10S4GyuVlytkMBrF
pusTmSVtj9P+am6Aqa1HUZhux13hZUk1BSNBEGPsKCZXOh6BBqqR7Ozbn4spoNctIfaz70xYsmGU
uX4gzNCNbGLWEM4ZxfS9t/LXeqsZoiZgKZ7NQHl4X+ZDHC0pbnNEIM2LIIJmCZtWEnKiZjCv8Rmf
tcrTwLEfdH1f0gZd7PXf+BiXZll+qz+Ht2Ngn9NqIZjMXjYl2LBmap1CVXU4kSR+F0sBf1W9yKNY
nUxS3x9B43XASUIAM0ZSQF2dhgA8QMag15agfMW6Q+IslNc6eqwrQ12us/h/Qfx74hz/xQ+e1JvD
djGw7WbwTQz0KdqUMhXudcc6MegC9IpRDOjeFlIKIw/p/YiSc/IvkxQb6CmJKRwZrhXp5Iu68HTT
2qovUsuIRzkQAAiXXddzAhrVjGdJ0siQ75c2VaW5NfAUcf6HNSr9WKIbDmjZ+x677OwV03ooSAIj
ZmXwaTup2TYZ7PbcGZhIOuH7HwbLRNama43bFl6tmtEo4PIgtsrWK2G4eBSuI3kzJZ8mgRaBuDBo
iR9EsFypDQMuKXv+5TyG9dhuMAVbyNTQ42za0lchr3P3236LGB2bt2aFsoag5m8JGXt/coz2xasT
As3LNZQIYwgpynIvmtacJ9gjG3MnfUGZG9zrGCdAnZVYbSUz6gS5KKotC2ScPAWkmsOYV/fcmeoF
0sDX0uwg6Tezt5rEjZMwEZb46DisP5raau9NJQ9W2+s8XrGnFUSEm5qIf/sqHMXX4sT9XXV+uV45
3Ul6qkptW+6aQ4YTTQZCjrww+AH44jfRpdSj7/rSE3SPYl+ywyo5Rjvqiy+lZV2qOzZ7mOwPP3LD
0r+f2mUezbW8hXjaf1z8Ew4blTHmhmIw5UZjEGO/ZYazZjwzpv741SKKzyiqtEkINPRQP0YFobfk
PWl0K7KFTkOFvO6xzgC0jVhQOphPA/n+8C6bR6oke2exSW6v6CeyVpweV6Dxt5QfEcRAb8q+RHu4
t8l1kFlBtWYj1qWe7sLxzkd5XEsQRiE0SwEB4INhj7EzAWciupB0eGoJUuCecrWUnFKT4khBV0eN
iFsZ/dV+ndMxBOMMtICqGt297UpI0x2dFsODxKKO7H+JXc1DGoGrtMHC44Y//hTrUDAv5ktauM+H
/RsWmO/uiUuXLLQ8YlMNNQe4Gbxokk6f6WX/2/tLabZMCgU8ee9Y5aI+K1xuWTprFg8ixzoEJy+V
JnmP4Qe66zWZ4TihtWGi3AMJPwR/wryUbdxx7+FNbs6QwA361Xt/c/lmU1nWptjfG73N//fecUaP
BKoWQdU00lpdfmT0xZMiATN1BMoe7+n7drKaKtT6Ccd5Tr8nke0uctwCA0gES8tsQwUNMENAM8Wj
bgNKHcQC85qLTiaF5AmkMl4v8tn+7bOnIRG7LA7S0ctVZJCdCBmKqTfpg8WtGnlEYgBGsvRxFR4F
AEGIs79cAjZM5Zbp6UuSKIYgA5N4elzm9oo2EALzaKpsOxU0o+MJ3XBrpHVo5I5VKKVK+Fxgn/JY
xrJdkGrGqxq8T9iXvAE9HBxWrzwWMvpNAHvDY5HDgjzPuWUuku8hSuFoHbzHjBh3a1G76i8HY8l6
zQDSBjlgPsxzS8f+NCN9QQtE1eL2PRKR9GM9VTc84EX0cAUEnpl6zB+iVpcuCMZqmFwoADTgK5lD
rmn1K35M9lCQGS3sYoeOdQy3GUIZ1MVTwLt/q7Zr/jy4MjBQL4fALA5nGet9lgVJA6akMi1JCCHT
hYTRWB2lJyWeNL2o1YlEmncgdQZqutamv8VX4ROvXmvhCNt1bu9HiE7+K0xVHZn7IF/ueMqlj+D2
xzlFg3Gb334ERLxbMI7/rhz9mvfv/Figd0nDcUaO1y2pXbqKqI16er5vWyHi+tle83dWMBPbFZb/
iKJY6M3eXDWUkZEAZjgbMcAV2Eob0f2k5mdeEWAjvSgj77ERG6R7Sb2qV1Mv9lZoCUt3qnJ5WUC4
Zkv7OzNzcgcGmP85r3/H9CeIpEgnQKwZwb7XSDYArN1eUK3+ITewv1k8mwgJ7jhWMgHJnOv53IPn
pDll2mh4wc42PnkIft0BOw0IMO/oEPKNs1zWq+dfowKCygk7NjpABsda2QriIf1pGELEAEk80fGW
l2DN4n8j4WlhBhtEUaxnDsvtsINM5xur63fpQELDIWhOe+FtQpOk0z4c6nAyKzWS4PsY1hCBBOuQ
qS6sY9sDNyfm8kM0y+Hc4RzfzqrF4J3GK+gFBdIw51GULRwlI9vH09pftnsUvLqodntBHdTHFWnk
wouroKLlfHntcKKW1YDPPo7gb/4PWjaHK8JamK48DWexbFiX9ddQtpiyyHVZE7GVsrDtHm5+BvVY
AhScEbNufrkpaYIsbwVLlbAIrlKpUt1qfDivVam4NWtobOecY+tFi8r9VBk9/Inte0yNYsFIweVw
+RxGQ7vORzXuJcoSoIFzzeUcnvtGOWmfha9QEhRRCHNnFDnU2N6Zaa4ELewsO1EXfGh5DFoTHkqn
XlKYb197r8nHRKkTv4+AgAhgIW+cnXpPxoJgJM64Yei4E8DhoExIeUHJsRzf/h5qbb5otriJSJyx
31/OMsXUJhTKllgcQhDJyPZiWuMabid9irkZyQPf7awmbB/DFUoaCwJBsZqMZJ5Fp/13LPcmaWeg
cGikhDKvaDe6w+DrBrDEL77xMuSyiUYsAlG2HnB+NqjHwNvdUlZfA5nIigb5ZLewwlg8EQQHdvAv
0e9DOgACK+ZJsMk942oGSKdhoya1b4dqXsJ9TrAo5m0qTw1dHBnFW080Zkx/gmMl3tXc87wmVjVF
oE/XsPa2K1SvYKYhLW5qwaNocwML76eLxXzXuMxacIS3VGKZbd7xgskF9qBSow8SzkqXAbvzYDx4
BLSwCtBsxk27WxWPb1UKnh9cJfrBA3NONVqTTW1Ql8cwOIgDoMj9yFIppOSVhA4UG5f9qu0tYL7Z
6dBEg80ysedOHh2J9tpNBJP5HJ/ubDR1tUAX2Py3o0DQOSrvrZbMxu6m1zOKMNu3RYJwid1+2P5Q
64qmC1LfqiUxBV1mCisN4TJNgare1LWo80CPZo5KF0uszmj39JIq/cgKjyuNbwU/AOUWnlbfxCib
Sa6+KYQHCnZoQrUNNw9Vi8XtKiijrGUotx1s6WHfOF/9tQ85V2QtCYPZwlyy51e85cdNucKRnfwd
jnQ4Ri1yEIznPm/hTuFNnkV9SXQBg7oeAR4d9ZRXJS28MvEo3qjKUaB2w/J0e+k/bjJoGvdKek4g
NBD/8MGme9qB7eXSVQf3X21A0NtpDhHnkDa39ySSN9wcLgCoIhvqHePNnlloXjMOOL3gKcWkLtiV
HL8xuUhdZ6elQ/UqYNDLv/KrlZFqrr8cUwuXoFAJbBKQfLuMKw01ty2LCZnS0GRBMJz9lFifQ7uy
zL7DNcPZyPGomH2rN7qOjDDAeWd0x9b5p+3Iw4UvSeriF2liPK1dHUQirv8AXy2LESm5Lq3/NLIl
/8jn7dOpTXSqaEtvxLtzGvQNomsheLsbJeyFSUE/HdwvX2wHiaU4pBa4r3fVjfsyhXIZuOr5/ZVO
xLpigG/Gzm4c14NAZVw4qAWLizIHqsKt+s9dG6xyXPmVaoolefdFLE/Ls37MRd+6vEP8T/cPU13r
t/rz0Y7QDt5T2DZJYx2CX2mOhRRbIXpBOeks7q5ak+nGa/VtJdg2IMUeOwdFnmoMTRiiSpBG5ZKQ
Nfm7uQfsaBGInHWdWbohHCjHAVtQaZWHBE0dU3stDI/ivNakvsJULDYY47cD3cL1Rts/BrTxoHLQ
MWU6bH9qARbV+ZJsQitI/HUdSdmZDv8RyJ6M7pfn5nSgEl4CI+oYfh4kqEQT6j1FtqjdyG8UnMVU
CHAFGrB/BZzSrWu/otllBLFYw1D4WTjiM1FC/xXo+cR5jekK9ywysmGZ/qN01fYp4Uf0ZK551PpO
BFxH2HqESaFgtfjV0ddcL5FPyIr/88HYy0Iew+J3tCppeCCV6XfEqgd90RSTdCw2p3vbVwAD49Cw
kJ9xaAlKHH9qq93Ma1u1rZBVjL4gOZR2cU46LUfdsveCgVaaK6ZpZqIjnxPLAlV7RCDJ+ia1H3Ga
dYX5DiqNuaRncV46QC3HSfEk7sLqW8yXXxfJ+AQynl4t6sXMY/pdZHJ+kf6j5lQ/yK5L7DPboOiZ
JHcbB/ogrBJKlzIzcqBQRru0H22n9uEMMAmh8Hh4ArDWaMZJrBg8IlPPn1bBIUIKwGNKvuhp6aNW
NdSGwatl8DZRvlH3QptWS4G2DwTDlAoVIUKHZQwSRf2br4UhdolItyPoJti9eykkEGYt7MFh3LZU
oWGGkb9NIKm1dGxasMfhqzZ38rvLDZfE3zo/gLNjNIDtdrrTPCVzqDLxhl82hmbF00eARiaEBCCV
IkOJNIXkhjM+cxNpe2y1ZDytGw/pqBd0frmRlEISRqsoNMZLbQW/8Xvnfjb0ezOwZUWVZY5OncXS
ZrGgKo4vU0j0Mf2uOA5z4VypuxjwniwW0x5DaZomKb65yZNPHWlGVepbLsiky3F2PEjlY29wKZ4l
5TY0XMhAFNJIzmcuLrE7qXuvnNM4LAU5rtCpVrmSMRuGny2BDH8ZjB3JQXjWfAEy7wvrQzDzEinh
hlKXhjtTS1xI8VoLpisxQ29mdESovSt1gWOaaBqGx4SWxgp4u/RDyl2sN98DBXgSFuNbHTwtRwDY
rbmPPB2aYYYnwOUafB/qgqaQ0D2m/9RMx+xUFAm99pfe5bruVENg8wjei2kvMREoF/EQjvmVfYkz
AowlR4aufK8FNxy99fr3mHoLULhh0i1EITA9pmcImLhPvTWpQMe9evnfZ1aWQXyo74W6efOpuGLp
g4gxhczj9Pz0pGsZfOuJtClsM4O7WmnjwvyZqq+Gj7fYcHylJY4pChvTOMvAZK+KYjp+e0ZqH2VJ
oJyyGIW4gaRGwVNc+Y+eAGoxHzsNND5DTV6cv6ynaFF72s3PUO02uLbsbg60ZNUZbuICR+K7cFbW
ACeY/ybOAKlz44M3TuLmS+opcn2yQp+XZ7ozdfz/P8vGKPG6AWAKm6i1K9Rx/xWvh4lCmrGI6b6+
8VL1z/mozBv8/GFINaqalx7bIUIDUGoat+FXHA3nwW+mCFpbDxKtBaUMrLbzaZWpaNSVTfIHmr3f
eStiq5BVyAQjdGbQEtpFUB8YAg0M+7tVK9VAnhjsiJFDBtg/a5B9OYZm8fyQoJbS2w8WsT4YmDO0
czdHXzqLe6ucSkJYWeDrPFsqZ/GFrjuPDDRe6mqlyKgRL2JXAlxpmJUCqET8cZTfVq8AKN04SDoR
jV1pQ5xs3c7TbiTCybE12RTSxvn8CqszYmPKcvMJB54oLxhcw+OcI1oqN1SynUMNirf9cBOQ2XRU
zC4+kd0X7FzRTLEWhvqKPJjgTXSvfvBerhArKLQAwSs+XogK1ZLHHX4+btWNT316HvqqvvTY30QH
IsULIs/WAN3t+lF7YnzXAMGcG2Bgn57K7v7SJ9WKihb1XNhnVWrena4/wE/MLyTOxzSZ8L+mZAHY
Yauwrr3IIw7t6yQ5cb+gTxdwbSuouMyYLPbi2AEhj4TOu57IbTavFSvuqe5SbmK+2ece+Mrg45E0
1FTLRCwP81YVxfqbzJMcYmQSwHbkMr2Hs8JvGP8gx+axrMC+YtPXhfB4+4OjF5RdQsGZ97VH0dLo
7rVx40CpQxjLNHL9N/JYf3bbaM0IRKsqpY3/gWwdRNAe4Sf0HA8La2i/JbScnhcRWG/9LO8cr1ok
SFTACavYOjTIo1nj/UJuU6gmJFzrLGTTkc/eAi35d9wLdFCu8br2PwPO0ZN17B6XfwR9/YX5xjY8
FhfVibqDWAcq/sGQhBdrIuqGoUPM5D9P8AfKZXp77+w05sbFf9R0EOzIY2FDqTfMb/OKcUMOOF6F
eTpjxEgnYG9wr1l9AHF7W3R1neRikMj60735yub7tSbNr/wa9BQ696UmWwDtxdsg6jSjtOLx057Q
OMbyxlOlg0uQw8A2en0vKRc2u5/E10Za7J6ShwSmJyRGjFn9ofYkclZkPZXScqDEKVEYfNkuN3rl
noWdLedqqS/P3h3M6Q89JuQRPMBi+9KZwrvHyuj38+5LxhRx0rkqNlOukjN+g/AK/zizhyZ2LpXb
aswZv+qEEd8C3NOf083E1LZ0MYV2+ZTHBfsGDNX5IjKvytpdCTtTpsdUuO1l4pejIlz4/iJ8CR5k
lJ8PG2sVXXPjYNdXL1sSiRaMHAijNXBxSBQRhcUtNdQv29o4jhsJHwYhN4IcNxTiGlxY/ebsHrqq
X+DQBqGr2Lg1i9c6XM/bEG28TNRuWMbqYgiGCepHKhOaQGQeZprCpFtMA9oRkzaFGYyEcZw2sntZ
N3FCfixVzRrLACaSJzrX+G9H09OGgjaH+EigaxhNnKTR8mXj9Z7Ov5xTCO+bwxV5YBaBL0gtFq7q
zdQZ7yMLHIdJHp1cVRDuP5BxSrVTCH00kxl85iUjvBEYpW69qsWA49nj/NyPOsf1dFJq6Njf9AhG
2fOtgIMc5Q5q8AsIjD1hGvk25Mqcb6seJL368pffxE3erC4A8Fu6E/n5aKw8lc9CDzQMECHVB1+g
JJNCMwgwdTagqXDMbqcvR42nn4rCq1nQeh0jkZraYTr0Key1R+JIwzizrREXDnFkbOYlZH6gp7se
FUEBe1iyy6XM0rocBlcRB9xyv4Ro2jJoEVKhhiqI+9fJSx8S3lvDfTkyGsCx4rOUPXUDlAo1M1Wv
kC9zjikPbW7Z+Rd/KgjTgMNJOy4vOh5UfA+Cnkc6SEzwVu9sQzC9c+DfIBDs9JUrHAIqBsOebG7p
YxqgWcejN96WlVS0a7SULCoTfSS71zvUnAvqA/dP59ZPMTljLW9vvrDTryjz/EIbuFetPpgSOcOp
co7XCvjZBMMwnsTkE3Elhe5Ikv9+zZgD8E349rFokKM2tFBlFcZko50OTzaQhS4vcLU9u/mbDOqf
mhgkEzHfI0mTzV8XEhz4d7BS+A4XsukNNNHXHKllplolBzyLAXcY3hQccq8umLGIxm9CqdRSNoVe
qqx7RiA+vI6etl1ARYNSOAedqiJJ1tSmmA8aEm2NI+vgdEIqSHhTzEG3A85L65MblXb141wRJcjV
Ui7O3P4MeTIyOe5yR1zLmXzpnoYNUMLmStiXi9nWFeVFoiyI4o4kvcb6A/XiyY7iXrktUSHdwNq2
G6QWFHEcHG7fD9AoaX4OToiKy8Rz8nxcPpzJNDpUZUsORIz+zh4sC7KIeniDV6sfQQ85eQjRpeUM
VDe9/zWCUStX5MY71KZcHHYPf4NrsLp+tsmMnii+6pUMgTO2Hm22URkD0a7dEWEMSR4BmdCI0T6d
3llXVEyXvlFYhyb+BxqcuFomBSHpu3QFjqxrBiQLPLlH4UTIWkp7uNrfvxGIKNXKIEFq2Qq1G0we
G8z8Jj0V9MAmSn+C84QXCR6fHsiuf+qVfeh2XwmPn2wb+nECpb/bzBOa59lYbhePJawlNtkNpnsv
8u3LENq8Mu4bIGoonCsY9ahmvZZASpfKOr9yTGpNEZf/kdqCHEuC2ZZY6UQ8EUKDshrZz9hQJUdZ
DXFRR8KtVJUplxevIsGJzEK2rQRZlsQjUT6XjBH3VEW0ifuVhpPqiTLqXkWgx2G58Ulq7+moGtpE
YfDlKUSa8xQBMkCsL0cwFpiXlVnVRNsLmE7IhBy2+ZOk7wSqEEzlUCuI/UDMpSn/1xZ79td5GNFq
SkbpjFgDTxM93+LTL7AwX9FTyuKMtHf4NRZ/AdbrV2X8Ju/6UvQVzhz2P2JvwNlkdDddtdNHBb/N
Q5Oq/p8vmteTApkO0fiz9UgbLW/veqEaOj2d3RSlCqzOnE1P0BBzQpAhq4Rj32GD//5/0VESVSLo
JpStDpRiJCMR56egSsPKrET/3L2igOImNaFz49DAxVgpkv4nA5k+okFZyyqpMR0EXGekjltwRfi4
wYEnbrvJreHpmEv+k3cQPNSH2uSXH3TVyxAnZB8n9bTwo9QkuEibEZGQHbhl9r5rE4zN1QL8kZxr
4GkIrYz2/5tccfIp8JqIAwVAxkLB3/WyvAVIGiJKWwX8RePuYMtVj7FpP5vG3Y5NKSUJi4ddIN3R
nzVCk/1Y1502GFD0VcjtnVQxLkkCPLbP+tfqXkehx3Z+EomG72DAUNrpuK1T5uuIAFd5y1AXpt8p
z1T/ArrGtUoNdRk4ZaMePWpYZiYr6FjWNu3igMWYX/+vkJ3QNqr2O6KqzU5YD3LaEU+CKz6auPnu
OpiaJZB9JZK0wvPRYkbpz+K1Uu11E0WKQ3NjdushrYjDhC56DPyDfuSNtbmoXF0xGezGNU+NdZZQ
itf0A2DzDy6ECYo8TOiv0PZHuj8m8UhmqYLXEI+3rGNdS5TXhe9K+ziN21oLAgKPmTpdmStmwI7U
0ieuvG7B/Uav7bsv6hCZhQhqlCOXYCk4vlnmx8TPwaaj0eEaZ5lhnjLoEykwYvfMVwBWBdYJ260/
XsbuVkMHLaiw7CQNV/F5lwIBk3eUEUX4i0eD/old6vNN4IyXSAFeiwt8+il5SwOjonxhopVHrfUw
Q4TY0r7+CDWNWlcXOubafbcnY4Q3fAUwht+wQ59anwyR7F+ktgtE8XR0GIgvJzyckLe5ydFceDua
7UArt/DgHqJFd0WaviO3rYockGfGJaaJwJHQrD/XMBmQmDE1pWjg0QvT1zlviS8vhn51U6eLpSqR
uOdK/cwYyTfdtNHFFD3iF2Eq6BP2lgjBOZ0Jvbz/JNftz8JMT5541hHUbPdcmNDl4r06ZjXKd3ya
eh8YOei7UH1/TfOV0MlW+DQsC7L4/DKlIWn7z/oXRCgqPJKo2PXvSNRCR09GmJrC0HAedofyzdK4
Wxpim5ZRoSc34CKDkrU2RPBvDYyGMNuJ6sRo1A3AtogW6DSQwOcdPlNcZkcMvPCfC6OVZRIHBPZL
BsP4wu/S2jgNvdAW3MNMeGWBqd97+qm0+sGtNWbfV4T/fdODXfEgSVOEZbGtf1EAI964L0dGIr0a
FvskQfbTPOTXOjpqxe54Iue9F3B5UA19x20ihb1PRgK8V7hYUkERIpowtulxLfx490iGFQCofLA1
sfvf140Eh9v7voVFZQOPLOLFFEgufYQ2s8Ank0BBVsBOuhtla3efKyDwoMayHlG8/asZ5Fkfjjv3
c+rzu8v2UavRzrE7sgqCq8ox+TsYm5u6SHn3lfeXauEjQDEJh88/IBl02CcsPSe2a0ldHR7hFjJN
T9G+Ppx4QYR57Kk63mvm9PzLb1s+WcRMxfWHLF0fXdqe64vNREPKR6Hb5/D4KvKzjrtlMlZXQCJ2
jTqHU1ZycMeCk6S1mI1j/B5QgQPecH8QVnYmPmQ3kDLVcNcDLDIYW5AElU7afhGrRcTKNIYfkbA0
8cqBhQhHG+DPeCNMJbHUUYRcUPqc36fybis2ibBTjTExilf+zgw6rRqhyBhnuN4NcF4kM2cxbl7S
408J5Ai9PWHln41qABsGznlCDbmjF7q3qMZoOUONfhKOSXuEquhZBpzy5LtXXGWyBBdWAknx8+Hm
YWa6fxrgcsQ7NqTSio1jMQsfd12ud9uaD+/hwmrGAV6SY/4LUK8vSOO1z2+G3110PEXYup+bIzwi
UWGN6YJu9ni7t/uo1CwyE/vaeYbXGhkRVXYOgRO43hrJopT0GmjK61/MqXHXeunozU3C5rTk9Q4K
JcvRA00synN90Ntd9SrpkMCsDx/S/aXFx+hSK3gsUtpWvdT3ThYrmVKg3tcuauNKMltk9X40K9zb
SgQrqOb43DlUgtcttHWMS1H5g2nbcWbsQL4biHKSTB03+nAu2EkFhWFxkFrngUE4mZGTxgps6fQ0
RvG5BGKfGp+F6/8V25reQ54iNiYTXjn9pU+iuIz0h1yhAC9JbbGWHiG9HZUan4HN2WJl+w7sI4YD
i9dD7pUvOjvV6XVgjByIkjDggjSJSStni+MPuv9b2G58JimDXF8xMLWMVEdc9Vfmh1bmaN8x2uXb
0RvMVh1yDJsym6CCiY+OU0xJhfCYrF6UwNwLIzm7Cr6g/5ME6iDhfi3SxJ57Wj2oiwV+1tlKLPlG
Eay7KHowvJ3BK0AMjoPFKTkRVZldzpjCPs3gcqrt6oKrna1usixaCP0vXZqG/jYugK3XFS8ypYd3
bG2gXwPY+WAh5LUKTJ/abDhcdXD/wVwNKygQLdpCwzsSyG/fLKPZmTFBK+CMBgozg/o0wINLTrN7
CmD4cHXbdATnIf19wFupJmkr1r2B7TRqZz9RQJBnXF1Of/lwf/EyW9bT/Soh85ty0p7Bp0x394q0
N+DqzWHJMfJdPjDGRaFRqg3hjzpOy7VCUnxgtg9ujZtWAH/Bf36mXKewvOHzCAkLXk/1Zw2bchox
FYwJscgoo+gJKP/f+v43IyZ8PNy0fVMYrSqCDGBUX3b24e5mreJvOhWpjwpEnfitQs8boB6nQP9K
3SZJbDDmz3ZtDjvARh55CUYLHnhskSOnXeCvaulD/IEhnXWEHff3tYTQQGfb0ITa8gC8AA3hX0L+
KvhfO3cIV9FnY5MPrH8jZIVVTn8aAQzSPx3RJckgYie0IM/G0atFJiGPKLvWi53jD+pFuY9teZEF
jf0mhWZAAbeqY1tho697w3I0434gFViGtH9pGGbKqN1F0TdYhf/tqlN6p5gybsYEJg/UiguITejD
Dmdsk+wD3Z9FCbLlNGO7Zt7OlJHIK/pH28xgC28Zve/ZvdD2rf/VaROe2zLspZy9FrWS3xw1hkwW
s6hIute88CkQc+ci8ShzIGVfJFaIRFEiweWVkuk2M99G9oDRrL/JKdBtbMIKJs51ek+4Mw3+Hr/U
r18ohlsMLY/KwoVuKCDuYhVdDNRVZE1hwzywgK9HVTKscfbaWdam9ZhNd2w89km14yjr6/N3c9cd
C3/ixbL7egE7hNneQS6ODKrVKLv4WQwxGq3s6DzOP5flhJJkJa24g3NfnXtOwfiitYgBsQdxOfaz
H7M0gcverZG3Kb9e0SRHxrL54Y0x1CldP/Rt45g0xu3urWZdbp5nbE7kJrGP6sh8eVdEpoYzW/un
ewaNc72xwLUoBEm3HI2MsQcAROj2LbLHTSe2TOdk/nr3qWBoKgrjU4RTlWMk6nxa2P++hzu6KT7W
1QRzEM6YxuJYrSETBWGbSq9wJwKKmms1tcNN6GLHFFXqjziyRtHMJgTqJ3lymk8cZSjk7K67BeY4
d7NlvsRSNjAwTQ==
`protect end_protected
