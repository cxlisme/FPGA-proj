`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OiQdtWTtR9UcO9P1itIuuwRl/QoCGJL59kbpJjiIH0R99OzTaBleFbU+NNejUoe719ezG39EaF6C
JkelkZJrEg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tfleOA5bEHRzyGZ1riApUseGRDF8C1zZETQ741VupG3H1r8eMsPvtNL8RVx5xP3cpYj8LXvKwLw5
0+FkmYCUB0nf19ebE4jV3pLqaaDpF6wA+Zh746oYvr13fHfYOjYKSPThx6QPXM5mV/5MBTR2MknE
Of/5cut58kXv4WQDH5k=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M6POsiNEQZUn8XpTzMUCVGZB3e4ppfCgsG9hiDQGif/W3u0k4dytULI+lkZzjwHgQak4GLxA9w9X
+UREx0EDd+SxWtFp22m0gypzAghoXKW7P8opjx47NLYnHrDCY6w5HhrJLdY8cJkwcBOz4OXprbw+
caQwLjRjMb5sTYBoAyuK3zPnh6dpAbq0pWjtz3eyNudpI42NkcRssLb1Iqdb05+7l/AK33vRTHaw
XOllspFzaXdakF+38oN+8uq0beSkI5kXfqakCLCmwvmPi7wKl8k8LNEJY+47fDj8vix49HTWOZS8
9ljmlXJYCiJT2O5pIOrUP1VlAIm6pcCn3HWB5w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dqO2wykDkPguKpl12j3EgkbUb61bN6zLFf7dCzJVoYaYvtcFi6H8lLOOzyjGJ3qdIdffHQNPTuiG
ssXPqvDurIxX36GKTwAwQW3ldInzY/1TXQ+o3jsy4hMPzM3ffkNtoljIy/lhMbFhiwTFJb163fD+
4HTzhQTM1GXIvyBGNJaq8GQSAYJXW6kOtUbM81zG9f+sBv5twJU9Jn7Jo0yRFodQlCHyKUDtTdPp
1nZf/pVhQQADfjVNYSJeV0pKP5dJ+UdXnjRL477weKhAFIaa8xVeLTYMW+zPqUGpiFO3sfAObidt
or9GredwqDJCvRcqeQI6xM+dIuFbHr2Dfm68nA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WU4nsMZg4YtntAgV6QkvPFMxWj4dZrhqRFX/kJKqJN7TNkPXDNA7Rhqx1+/6uFwuSaI0AQrdxFXP
EVraYBkDO0RHDESoD4kwhhn8GN9o/NL3N139r3nkl/uXc1mgsluDRE/5xRkuEs1iqhdeReBjBBh8
nZAR8dpdZ8jyt+ArMP09QeO8SiHiHRaKjEhJj1pok7j24ZZjJYvbmJsepiHVEa/aBvCK3h3JK2Fk
A6kyTBcSUgAB5RxbX38w7XuR3X/tG5FaP2RdqxrwN86cSZgpDAs4Hqvh5h+F3Oe2i6NVVxBeRsu9
PpDzdIZDOqiKVW1xv8K1oGmvMF5aObJ2ctzmVA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FyB17WZbhJVBrhgthXdKrkqOlqvFFDagDfs3WivMvudkE/iPtXeE0qdpXYAwxYqNoWDs+ElK0mAO
2kolOuBbx0X98agvv5awOMlh4eRz02zql+1KckZ2kLYv8NccdLWfYupLFCW/JSgJoAncjrm9qrw+
UCKXIVlXucr5POaBUpY=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
s3atYiAAjOvqgT9M5QG6BW4Pgy2gbkhbIa7BRi47fe15EzjIBPGwNinWEHGfCCH3/mBvgHwXQe5O
Vvj3hSf/mN4mHhJQVwCuMPhKJzTBztkeAjcRZaphRf66A0TNfWY+Xt2x17GEgNN331eisXF7v9C4
5ZUgJDe3v1TWAa8ZmTjbDhgfQXsPeZ4NuAcomX0zRSBCeuwXWUcDJR66TOhpbpdKVRa1oO4j7xpC
SqtGZEjqFbQ5kCXxI6375ZpmuyI1lmIA4tSGuRlC5HehcCC7zoasyR9u96M17hdwFJF6dOu8QR7L
J7FP8imei0wQr7KAis6WAmXyD6+ZwQApEKEcMA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 60560)
`protect data_block
ntlD7e+Q9JYZjDVVLQFFcmdd8FyFON54X7kspq6ShCefmhLBaoJnMRfyNlCgh6+hrb0jEk+A+i4W
pdSarNyVijpiyRV9Aw3gA1Yd5gd6YDTdoYlJxpP84i6Ts0gmLfJb15IDjRwviSzuDC31migiM5dE
4KiJJdu+yCpLNTx1SzXOWS5cj2IICmdoA+zXMNFwwnV9Qia5O3klJE21xXNPplkOPGxZaImJGqeX
bp7IE15MpRZzda6PhX5+OJDVpROl/Mmej/lAaH/6gPQw4CSwJb9Yhb1HGygRUJsQEf6wlw9XkTyv
El1UFV3YW/TcC3m8aCAkS6QvC4UNRHE/QsfZFGWA55NrFCiYaRqB6BlqgUCrNYh5cTQsWiRGU6sY
/ll5vtwVLTqMvc9LA3P02cB6NJOq7hEh7tIgHmNarnrTU4kS+B6n4YwjsJZY09o+KD88tf3SxKWo
UWpYYUn4wnNb7xwD5xhGLSLK3dF3aYo9k5FZ7oYGJIFE1nfy7s++y6zAzFbGHhJHdPPTk53oFt25
qhwLUs9zC9HihTMyolmRcJrBWegaRdc4aySo7VQGIwzHFGiQ9VxFl3jf7mSgiD9dpEb6gsWEmSTG
1dF2OCtQPviVmPDCeXeFcIFi25ZgzifcFxHwbPEg6AJ+UmX7nYKKdSa+4NAhJw3z2c+9HwZifkq4
5jmMr49aSis0DpBvuyWabeWpj9zc75Rc6X+y1al7T/h4N+3CTUon8xe9s8TlQ5ozjYE1t3oIH1Aw
gJxIzp9htgUiu/aTpbiAF5Z1STXs7DSNkTWbVjbzOO3AOH5M2HdmV/Kop1WEcb9quG3S9XEN1TSC
/A1stYrhUWkS165KfBTEIWn6CdYefgmhE3SvqoPG8jgJteEmwkYowaN/doyNDMwZO/J1n6ZPe+Yk
4n6uAxfFUxla7cpXoIsmcGmpiS6z8cr3opamIA2MBmeLfzHPrQsKrbgdrd2WItWDcUvdyxhOviwN
JawWLrWqewzK+o14mBDn7o4Cd2HqbRXfSHZqX1tZxTSQDwB6W4AKptcaO9HH8E9X5HeZTlCRMpr9
xPMd6X9Fbs2pKy4Ns9vNVPhhdvybOzGFn/W1j8prr+yvMU1RnhIhnifp0ziwYnHTJQfEyjAQu9JT
MQQ/4eGiJR7rClT7Z60iHYrRhtVQ91T/zzRgByWhUYIpikiHPZjrcuuB5SPpeatciYbhwI91PVPD
JdkFliPKA44OT7Z9ZuIN9J3CsBYbnSQFMc3vJY5Qfh41nVSF7hOntizwtXGRreYx37mT28mxQJg7
/vS3EGS9Q/xbKMJRjiKwrrOBWj5681YTqlAlVa/9bK5ovjAbd4f1eXe5ZTmuFTZ5ntYMiMic17Pc
QdVuDR65AjS/5NvzU8lUgeJCqDTNh/wi2+Veb2veyF1i6GkYcyBSzngE1cmbKbm8ArhufADsS6eo
bSdMpygKCA0wSARojmPRVfAvw0dgJWvI/nO++/ATm+S6WqzW8CAC80GCz3HoiYg/yKAfCcJdCq+U
lBmx7UDm/PRBNo+8k7UvkysZg0pEcdpQoQT5hUavHJ3ej2SR9gc0lUQP3WLRCoPiV7R5Z0PPfCdR
5wrmKJEl1kcPoM3wbud8e9am5OouvTm+t1KCbHrDBV+KqJ1h4ccjNW/JrNJSa3mb+iPueUUCNY3t
JfHZnybbPQ6c6hMtiH56gBxFms7rJzsPGoizcScoufEGHslJk2eJf4R4sxxwtk3jNsQYeCo7oc1P
q4tlU4blqd4ezLZpMlbZzazjmb/zx3IT6xGPNcuSBrVWhlPLBA642lB+rxujyGn7opn8DiElwM2z
FxNByYCymQJSqerWBXGdUGUK4mqARAyiqaQg+uS+QH+fMDrm0uUpeRPTJm6rN6/zXjGuOeSQ+VS9
k4to+Ay0YuoJAZGETQHiyo0/klvjBX4ggVYtk0YRtjrrpaBonYbY00R6y4XMsWtlcQf7RZjYskVj
0Ks//kreX/Qmo0iW93Zr+BZ9P0iszvDWvpJjdXU8usPkP+DySRVjQXNGPv5BQQP0LlN7c6mgWRpW
fBBFTrPdv6JUov99oln0GF40LFaBqLvDZ887O4oW1OWNnm10eqYWUePrgQmZlzyt20+2c+3zLdh4
xA+os0q94jZZbaVR63w/L8N2BB/Ia5QRuRX8AuWbvq1+awghJBAqQIYKQaZJiGK1tOm+JzQOfuPb
YzjRrxnBQaIZb1rnj4dDwpU/tJ3Mk+f0PxJ0NjAV5tPlf1GRBjzHgkK+o9i1kwNTW8wAh0u6UPu/
leNbmCfUr7LkIt6HvD+Lad+b3QTGhnoYm6gSGD3rR+I5r8Hwxrrta2DdgSfOM19j/FQTOJgz+MkD
jsKn7mfBvMP9TGHser78iKjBGRofkyLbiBwvpGpl1qkN+lQSCef7ryVDwZmZoWw9fdlsvoUNukCb
eRzXmMDD8rw50v6NoRrHjqHYQQAmvSqG4hkGCVlMdh7JfN/QUBiEu24+kI+vA+ZKcEfL92HTJGrq
bgOY97akKqa+e0olUbAWM6Rn4icaL/ZHiR7ep4SPYLysbGBHgpK5tUA482JO9yghBJpVcuecMMkL
zuZVdDYo+Ug6lGAYS8HgpfUg1ek4U6pJSLAMDxWr55YeFeWBrV5tVqeLjy9WjEaMb12RSC+HAHnD
/eb9+o56d7xNWXr2QIo1cluAcvsPKIO+asQ6aZX1KSBS0L5sPOAvPuTdGsbxY3fqXlOT9K8XApon
WlkDckjLKmBb5ARMOnk5I4ihO/qW3nSPisHcPx98XZKoeewjJEuIY+jmwxa9CDlkoDKvaqT6/NR0
vncMzv03Fb8jQZzzOGC66qMuXwrYPlqNDIBdZV0HVpgG3SUTf+jnKIiWzWu6LtYHjubzhpc6/7xW
aHrkl2291uxthib1M3iDee0mhmqmdf8BjBMdqPa+vVRVyyZTWiYjhGiIeK/v8ISa1N/n6htDDP2X
p1dbhQ9WvOvYGnLabT5hZ46u2z6wff4RKQQsFznizRBpXRGex1rfwrno96r+V8Vd4ZwJOU2Hj/vY
zEORl/xOmMNTONjU4BuvLBU6QzUNBjeEPsmbC5KJ9ZVGMVFVkxZRuQ6Vn0PW+KjdG+xZZkN12YV2
6Q/mjyatwK9k7yEJjAXP8ILv3vXwMVEgQeeNhpAQoluC5pwuu+3ZLEAvDdlMTf5aCqUnPRN8BPJf
35p7AkMoQCU3tWnU43EqWOHL55i2+T9PVDA//IZodM88QivieuVOwF+7YJuv9bk86Cqsd4EIZwUf
yLECRbXFzWeso0UHZO0qT+03+FqNZs1IvwjnvkjVmB6T7NKBv27qJn+U6D0NvbKG8UMuWLdUKDzF
Zgl5iLcqfYbFL2TgFeCV6b0z9pMcqiPM+Q+CnmLeGZX2LZA5PxQlnlCyvsORxx//RXDOjbZRXmM1
sk5bYUSEgRYkLVf82OTFXKo9SSeFGkpyeIvxRVWWt8ICsksiu25FwaktsnYGRPGjBdxopRmqrw3i
wq2bv3Jy5Adenf+fk83eC0H80jj1mUbLNbnPrygASu3kA3lmi52TOTksdmqzi9YzmqPxhVf5QY1P
OmD9XB4OBhbogOMEMEwfI+FKdCldciuvVo+7P9aYSIRpKkCJG3oRyhLYspfyWjgS1gvsBIsO6kUU
ZX6KRmU5Kc8U+QEZ/o1pRqpji19xMJPflxgK553oUb+DTGRiS0/bb/qH9Ef+PXIVqMX1L36GHnHE
0DnUuMl6R9sEJVllxrZ44P+7IJIbnDBHZnMKxX4wnMY17L2ex2iCdvs7wLFXpxZCmL1vJHO1+sfn
mVHIiQpTkLB8DswiBrXkO8rcIJ6i7u6sBQZsX3p5VqUerQUAV14rh7R2bNgX3DYiuMhYcbS8oey1
p27qrXWRwpgFMlQV9uls3yIRNWl9XLep4iP6qbrHgZTVE3jXxH/gx5zip7GCyRHmDpLZRPMOYVUy
KATCTGmGd2SSaqIQQXvlFLECBHO+8AQ18mM9Jp0mm5rcdMv1PJu/bVqepU+3AgisR/4bQOrPxRFQ
8wbTI02EhEOQV0wr64nO9JQ4xhsbzriz74TbHWZejVspc05NO/cettC2H8dQj66eRxYfAqV17mVT
Dv8RSWEZhseZMSPt+fnxn7K9l8QXlHmJzsQNMKdkya8ZUlZTvHV7Jze3/mFb/+WBAq15rqtZt+4o
TCYq5K2OrD7QuSewGfB17SOc5GueOP97NV2uJvQsOUiUSXt4yRQG7UbSM0KuqmjZBpDXxMmXUDPM
Ql+40YJdTp2phsXFU+GBclDjxFfVVSlZ+G8+BasHo+EFtsXZl3S4ZMRmBE0QGDhKznKrIpWm3YXW
R1Cp5a2U3lMMWVJwdUeml3gG/vN0wwE1nSUTSMZbgM1Q5sKKEpad43MhtkZN3ETSlEqCWwXk/e7f
C3vAxFkVRuYVdRiuO4Bwq4yAcmwB0lRhlSwnb6zv5Y0isJ4L50zcj/L3pPbAlA9PDa6gwVgUPLFU
y39kiWmL2uV6DPEmC3hBb5rdqtNObIicTFUasepqCxbaFjOdlyFThH2tLI07Z2RtkxEjeg7Gtfkv
80joLN6Vf7c4UkBbX9POptAGqXhx0fL3vEEqsJet6gd21I4+odXTlpHUD7SKec2iiSbidTeFh9SV
NySR8OVGDgJBR2OTco42sNhRjZhpqtzk/7yOi0L6zyJySZpzFdfNdhcPEugwjqSCWUaPnYfWkmRL
77LtL7mh64clA2luqkwoB2+znPDVSas+GHzGSLz+IdgcXl3ZhqwIDV8RvGqj1ct2DTaHnmzjnJvt
kNqe7w0fQ3qPeBClompf063KT+08ul/+DniysG60WT9RHQ2UM5OtC23rrN518D8HuCvQBfiUno3R
JjKXQYrBF3WZc9BuopWW32oCFePgXrOwzfTXQAmD5l/UBwM+J/BELBhazUxftyMRf9IMMaemXTqX
yEwtdGuKL0flaYs7t+3n14wHXZYZ7XK2G/H/+wJajqQyN9gLFiJ9xvFxzAXayewRD/EgrgjFaNQ4
wb6c26yCqLIQiDErBV3BnjwhiFjWcpEoxxmG6o5ImL7APF6eBQSxzmxO3xSfIiHGKuya2QEBRXkl
GNfcxuXiQ0BU8vEB7C/ojMPWrdkBa8Sa7HIe10vrz/Fa/9qqYV9K0Bxrv14xBC+WblINdDPyb9e6
BoAnmCPC7PV2p8sBFwKek2upqTTlWMZ32pxfu5CPFDM5wPbEPJnqzS224ep2nQZlSyZ38kZNhttM
JMgCLu6JzyxYt7ZO51JNTffgmObKWQPiO++ldVQZTWufjc/o7VTfnRMraq3h3Fdvs2mCwWi3HUeB
jdceLu6c3Xt16OEhkucyuMiOIAREuXgb8auPqTToyltOYrM4UqITUYhvKilaIkoirErFltiZ639S
NhRzfmLEDFGXDysI9tGI400m5REo902nOlOXQQRlNZe1OXcYJJtRYsSrKc/j6g4gfhuojV09iZsS
FpTv7WZ8GUbNxb0J8AwJqxYftzN4HJfgv4LuV6fu/3epN8q0uQBOHH3CBNaYyErSjWgUgTQJIgat
Yc9l9OiE8Pq6C6qNXhBEwbD4o0vWlJVLVKlsRdwJflAkKCWDZsD7rCOnKRL6NjjnYyIP0jRgQYgN
RSuK6F2dygL4hLKaTdKaA9kPeDGyAB0AlJ3kSZ6b5l5R8xIQlbJW2YkNdwvI2EAUwYll/R8bgKrG
TfUQ1U+9WmjF4OILy/fqYlFrfiMil7Y7BUpSbOnUqFx0booMLRX0IjuQzONbJVcSmxOPfbgvTF3v
UThls5oR4yoHOlmAscwjuREY1+nfkFviZcxYHkbkrXQN20ub1ozTnboyB/0OAUFfn2LWVnE+9DW8
sVBcEm2gFkSO9iDwM2FuesStOkm69DqWwxg9s5aYI4d7ZzHSf+6eUZBav0xpumgZmwoSup98w06k
62zYQ1A4j3kOftIYkYSNouF1VP7Ch2cwL8b1t8153JoEUGHJWSrhT1cxgzf30oBZlP4FgzQiVESr
s50/D0AFIC6rMK82IyhKDg9yjCoH48SVcaJTL4OltNL2EC4JtqgfqB3yq6ouO+GSdB+MlM6+raDD
B8pZ+z1aOsTEd3UWm7PI7MS2M1hn1Q49+u7zU6V+1IGqSJEd6ZT/s4iaY2+07D6yd0ThkdnfQtVu
aQhscrfthiTeglcEwD7a2jnlr6/VyvK8TYhrT1l9+E5oB68ICWrqXLefZSb9ETaEsIQqU+GVNSnK
xAysTxxvFisx80FnMy0MRBSwuiH9knZP8bixH+mlUbx1RfKpghSxVlcm3/UjqQs+vGpLIlkn2m9/
X4W/fU19Y2XtHN496K1ZvdCUlSxzPqRgjfiiYGvvikArmPmSmBC63Xd6X2j3JFWSHncV0qNqj/C+
L+GRZt+v6ozyh/6Lb56BQg3XmgKXtJLDBYrd9vmbNooVo9aQuiqPOdNa5xKGVN8cgZ2QpWI69JXw
Z/z43IEWMqs8MAGNHKvU74GxZVqYy0MET1pJlT0tpgz6RzsRC/ud0HymVwKbPUzZ5K8qDZUXMWtq
60XTxvdSyLH5APA0gn3syXCVm9me0z1zqMaHh57cppMNnHeYVaBLnP2M/V+oFVnR0X4VMITPa0li
AHKAcaXmXkU5wFSqMKJnODGijlkWUEoUeBOPH65vWsn0AaqxtQ4+0eUm8erNLWB1AEt9AKI7VlJ3
8bpMD7mm/Fhr2k3y6GGgsFLjqvvnNhnOyXrpsM9xmWfTGx0Sb/sc3PEWEu+KNvIX3/WpZCuHmddA
xTVHT2CAsSIwPMt61BDSFQjuQpTGVanQSVGYl+rFkDV4kRKPIAaKDTpJ744TlIMqePyhWg0rQWH3
bLmW/gZMTDjKrg7M39W9DkEcRGsAdNfOg3gzV6z1beVvIaU4SQBTQ9CvwkGnnFZX7wurjqMr7xqz
hBChiT7uLsWu7Oy6wKLwLprZ6y5FVKgIQ43+DZ7mRNt6mJw8A91ZJGNZQ1SSu9LAGpCeeOJfdnfk
X6Andz8zgNlWtb8DaDLRGkqnpAOKOy7M4hMb0pHdrTovzMsLcWDSw1aJDEaRmSoIRROUuouNBDm9
gheGVLDbbPCXBtx3CINEc1e00uiUpZ0P1WnKdJBbTLGd173cMzkbWnYgZ1lisZOPGw3A+y1N50jc
w6Qd2p1xXSV/PdmODtDSub+l2GSIfMiv2E08Q7sCXUkEFY/6d+dk/BJvRFdBVDlxo0jHYvNT67bf
23+MN53d+eHYSTK+NQ7FY51kpqXMkGq6Q34wWGy3+HDDDTLeb2XHcNRUmwfo37TQcdXQAJQLHLIe
l/zUgLVs/lKM2hc70ZBu7SJnq4QS8ctuA404BNdpvEaI/QYQG3J5URk6jMP+NHFWVoDUVUxWEXf7
42p3Irzhle7Eq1hg96xK5+XJr8034KI5ycGF5onjW0CDp8QecjbCCsXiPij1pQjKyEB5OrcNCTdm
E8gr9D+1fRXV6NcS3jhurK+FSQGNMSL3IIDjIb6EE4jfgw0VAcztCOiSAexKDjIWRaXfLrhMDTrp
IF/BpgOuR/U4jKoc8V4ynpJuBqcy5P6WVDC3A1XVS/hQDc0fvYK7HqsclIzsmc84X5yqUi3IfyqF
XuuwiJswsACpzXOYGPFRQ4ZXd6CMV0ZvAizzH+cPTp4cskgG1OGBGfh7yhcaPlkiX6uieqfmkFVr
TZPlEFHeYnhFOaB+GOpT8P4vu0j0j/On8J/jkt7W1lwpTxcWrNwBfRKL7FjZ4Ai+YWTakNfe2Svi
53b3X5ukqFJvIDQ8Z6wwCUET80gIHYfBgpVEBuTf3HA4g9QUCOjJyqfG8aagUZ7MNIAliKzOvH4T
g29SYvmK3NOLMsk4jnRcBIGIPgtD+AGHIEkC2eXCEegHF1FTTfuw5wnmAkZi+BuGuiTlDCOoKD3T
dpsmOxlAY6bWhwAhCi3ByAa8u86g7U2T7cJDlZsy05zoBV+ZbsDUtIV36dY00k/xFTBd62qRSFz/
HxBgDOFT/s5Tl2WETNmVQOt0cGMCUBADVZKRU0tVZp+3LHAZRvK1BYlCVOmz+GfUFxNh1E01+wFV
uruYkZvuSsRU2oz4rXDuOFm9L9j9Z7mvoRuzSkJkdVU1XdqVtShrgXRIcOJvKlXT5hKOiQpSGYAf
z0R1D4mYy/+wMUBXM3Ol19fnNcthk0Gh+tpaYHFdISM0MJuYGINtdjmn+wTLuaiP6Xo7CCC/SVIO
T8bkzHHXcHHasgtkcma8CtECdrV221syz+LJRTCa4juC9qFsn5mmD3GTz0ey1iTbUcwoMMNZXMwc
ouICF1HZJI25ZSLezK+9dFD4tJ0PS+lm6D0ZNmLRdcZW3wLWqUYXYQbOfQ8LqrOnLKodqhigdieN
afuLT84Fa2MSoJHa3iy8PyqTHEpL0U+v3g9AnrppbEAmN5a2gYF/zF4QUZsA2pisMLjaDYKAPOyU
e6PTWklnUmlQUo+znt8SUlcgAXwo8w+8XD+7MJH8n/QPixOFySVeSTFrg44ptfcILL+sqx5glFda
i2hVexoSrDNQGey7rpoP1z5pnZCAc/ktGbyDKrwALU3MKrm9qY4XmRoFuqKL1AfV23Vunr5lF6Wo
BB6YBNhYB4lgDaRURp3d5bAcsARv/i2ha1ufDRiSeYIB0DVUHcZiwr84cdAaTmfOhPFMST5RGwhE
DRk2V3q9e5HPdKfJZcahjnSPXtFa3do4lvGPcgIDhTdrwQ7QtLCLoGtCEPrhrrws1gBZmVju1iqr
Ctr0MONxzNb5o6UY1ISbjVQaiKj4APrhn8vSv5JNzcIqFmVotC7ac3mlz+8DI+zjjka7VpKFQePa
o6hkVtySBAxxlsBMdG78DbIxRoWOhk4+ME0ckMDE2BFe1O6aX1D86wkxLJkqV2z5aWAlxNJqk1mg
K05secMvkbjPfQxsxYx7lV1WauFf744YELeikP3UETWcleLLvPJOFMWHpG8K2pehFe6tKsPbJanY
cStEUSzGkZgQdmus58nDZ8EpX+76g7t5IDryDLuK06HHNB6aIOv5jSg6v7/NR+yA6LghKpIFUJxi
UkCmw6hur+b9ggAHwaxbTq+Igmz+ezCkAevcQDxW3YS8Q4GG24hWKSwFzc35YIoV6XPiE8Ujs0id
ax4tgnGQwUI2A4ZT15MoSls0fEgr1kb66HaE+2IaLw+dRslh6uOlqiwWf1dVyNFP32LmrPSwi76I
H97Akq/Vi5fxX3mXmVYqlhQrEYtXy9U1/t1ZhpnlRpQMcwVmLabBk5gU24YutEF68UTSkEjGfakH
s+qrps6cDxom4I63w2CSabtLTTKBNMOagWHty+dvHBJLXh1C27mINQ4zOmIvQZgw0+UjKOZNTPEO
aPjwJXZ107/pB61TUT4FNksszMS59bxRxbCJafSczbdK+j1w7DZsjyXH+mFnLPhuGCGhceqL2qBG
8hlMIU5Yty2t/QzPpYU2+MpnuPIsr9spomkFvdd33Iv6krApmUsZWwdi14hlklYWVOCqkkteidrW
JSPxlk9BPsypgW77IjQrLnRbU2dQ89zg5watcgNE0zssuFLGhGUpzydD9UiLNvHVruu5lsEPuOHn
fLJyaN38Vaj/+VichFWsVHIP/dp6GOdUXOaXAgVC39ukwZZh3bt50WSQeaNKDclE4cO3dgXATQZ+
CYlSaWGT2b1C+9f4Q4pjTCqbye8I0gZ2ZZV80SgSibmWF8FHWb4zo+b8PUjdIkRK9ckGbQjPFEGs
3oNqBxR2CZf7h4Zkw7xAdW2zCSHgAFw8AzvOjgbnOz0AFhUKAnfmVobK2Awwa549e+toUMSSwY3i
SSZ1NxfpPzzLjgT1ZeLY7nV9NDpB5W/39SzLUX4rkMuYKPaQCaT1nyVXESOT3AJbXqpq0IF5g310
+0QzD8QX0ATQ6K1NihTCQHyoowhNKfh5GjnRRKcqZ2foeJE0v2Y7P/4xFhAtjChWyCuD/gNsnnDY
qgrS4kJKxT2+N8Z2VbtbYhxRMg3inbknD339yGJABu5L46xAHCk87e1p5P0yWpoEL8djHkZOuRSL
MWx8b3YREWA27oct4mZtKd6vK4ORuEoOB71do8o14YxcO/t8gcYAyFNkG9CKCIytHjdIHdwEqD01
MUfa3aeu1cKH6k41N49Cf3IjrdmWYEwtRuvZaE0moN+ZSFYNoqLZDurBF7kFSpAOj0plq3BglvUp
QNZS8Ajm4eDuRs7QXrMIftpUgiwdOv1wlyDBJwzaAmprTGLI2q9yE/cgEBnvWFSMbxV34N6ySxAT
MWcHrLRrcOqLgfg/b55FYpnhy32vFl+Oo5inK1UW652rBDuuf9U1JOLpwpnyDZX7aTXTk6wcGN8Q
hcwORHPrtvxf4OFer+KmGJQhXlXlxLKhOfdoFkHKUgkr/FNgNkePK8jpKb240gelwVwRWodwEwe3
Bjh/AHcM5hKMiNXFAfJ6afMtnfbv4hy2ilxnDB8N64jl/3NHP4uB46hBOK17i8iuZb9qfDh1TTMh
2a6Jiy9D0Z+JEHcP8N5cN+cCLLBnFPoLM6CkZzJP2B9piJDjSjgiUQQ2LSsnszVd0g3Hx9eBTWl2
bQQVJ3ueTYe1UBQqaCxh+seJ46Z7gIkeVSBw4UIQib24ixwp1dSBWxy/on6xgr6UsZeF0OcQGW5h
GoCW/O0bFHiM/qBPX2GvcUhzXInaitfetrTYqZe0jBvZFmlofrVoqwazkfK4ovJSgebboXmj17rk
3gKpwBg20iMK4wxBb1w+DZpVZuFqTzkbs7BdLYc9mtbZKKnTW/mdiWpC3eNgf/PD4CQ81VIibdy9
hkRko3MoKSPx+sFpOG0HmudtTegc0XAs1Eds7NTyU8jCPMk30bCTYgPHEz9ujz2eAirBfL8LC3aY
S7JIWK12i4Ipf7WD56FnNtEa7QYfethirrQsAzKlgEIVvqNnxN8lvGqfinT58PLkQ29I99JAmgQb
9t0G/WfzCAOKloJqDimUO9KDZEO2q1Ff3HMlENBzD9Py6TpzZRmm81qW0tK5QxP1gB+iKkTovEp5
1xyFogNhQPKCnnVcZwfQ9Nm8SH0xVNuz0imtwT71B6B8lMMVac3mACC8vc4BXqpUhFhpAOBvifyF
UXmvPk7YXQUEbFbqJD1FUvkFOtx1CQox0NqWGeufPWriNQrcEG2V/V3D6BqC4XlGmV7eBY60k4Pr
/AClh9o4WaiHYCqLVFB1sacavWcmDWHlNkcIx90dFLm1DN9mqteMLllXxHGDc4Tc4xu2TBW4XFJp
l10Y7ruzHsQWgC9lsTQu+O1kJtQ1ujt0sxVD/iP7WkooZfg5KwZp40aeKIDOrTEQnW1470bTfENK
0A8c90buAbfSVZFKCE5vxmUirLv3MD2eeOCRkWrpgfWN3J8RA4tC9FvelXN8WMS5T2MMPJurG2sC
7p86oHzP6u+L0AZLlaPDASpjQHminUN++/WJI6aVTKotgrXFxsAC7UqD+GEhnTugSxKUVJ36q4GM
TQpzMLxiFfo40BgnwZNkIINW1MNPhNbo5qNf9WHNizoEQSDXI2PvigIjM/6bh3YiBfk8w7gHZvEl
2aNBm6yEsQFsiqofP97PbJ8LwyK1QUl+h+DzhMU9v3d7h1X28KhZ7vtqmrktoic270t0V/JpnsnP
qwFJ46vdWPyTpkyxooIEYLV9USZoEP+CkMLjk0LQPolpUv/IPi38d0e9rotqopFWMt95cYaWtNVY
NpDfF8y2kYjI/eycXhsm/maXJBEWntnW+wQOBJ4+s17PBokXEkoA+29zQuEmtRfvdebz3Oy/Iw++
WdR2j+wcwyb6TRxRp8NjLFh+LUFByIz2Zi3jC22iAnuU6lCjoIMU7fBJ1ptiIpF84xao2XpgwZGc
UIVup0hr9JW3N5XBIfcoQv0cxRxu9jQlOOR5UjzmXa66AZT/6aeSL9YU20MXSd58buSF1PU9o8jz
mG4IjxjHDNflFQ/5dokYEnItIwASzKyFuX8DD5HC97SjmJ1Mt7WN5hI/tYkWVzLGVLm+pKbN9a34
COJAkjtrl9WHUcAjlEfcagtt2QH9KoObASyFQGRWcpdWbXEKA21DXC08b4NqFqTVdxfM1mj4c6go
ojdBMl/XOVbBsNRcSLhe3+OXC6p1MDQ9Xqj6nEMGBfoyD1gYt0mms4dKZOxJQxYHOYHAtGcM5gKT
o03tKHFxdorJvEycM6qNZQjG7h6djKNiK8pL0d9fti/kmWrmLqH7WsnNMF2gZ3UBPuNmivLCqQ6s
340HRNiphalmQI8TMo03DWLB1BMDzyCKbZIto0+qMw2S36QrqINMulPMyyCPwf1VXEOcXyC9feCj
o6If6s+4QGuCGcFYYvm/+dk2FPOX9sND2q/mJ654NQoCxax2W56MrsPaHjYqze/JmC9JldjOzffk
LLm88qOVYYQm3MFWheBvFp6VCQIGRPkm20dy9F4/u3RNWq4GbrAddFX38mJeSMvkD9tKfg2GgCEi
gZig9KUzTRnE2qGIBw0dPEfwUC5Bl7qRzS2VsTnI43q2BWeQ1ns8uy6gBBMMoPcLYFAggE5hOMzl
ATv2SqRQ89XLcVMjXxXjrxw6S/5cPbJOY6AHDOVFekpq+t9UaE1V46NQw7SqUa+zNthF2EEMRhyC
n5rZne5Rtge9AIel/fJzJn++gt/Wyxx1k8/6pQN0onOLzybjZZWj6P/3CsQYapLyKXawPSYBYTLs
7N8UvuNtPIrkLPZKF3KYjWysQT5n1LcGmFBpgsJLhdT2R2qrcYUqaCMrLGweTs8JXvGX5e2rWAoa
tGEPzCRa7eQ4UWc9TuLmqgKRYPtObBPm8J4R8qoXvmhQEXvpjURFeRbAg182QbYNvyqCvMAmQ5to
RPtfUSLcduxpC4seOTP8BYKnpH87zh4jfrFOeKp08YTFHSwX2uYrxYoCQ3/eAzbV2AROpT/EzwMm
tjBISkGZ+qdGr+/8qBoxPecJ8kCF7nOMtrS75DGbxtrY5RO6cmVoKjiDtDlPbNOoz5QaGrUw/DAH
fE8/pxTTrnY2ZjxbnkIHf95i9juLY2IF1DdufAZC12K48S2O6U1dYttd+/9KL7E/cD1STWOKy6XO
fh4dFYVnh3bzZhcxV+pOLSApBjugxBU0weexfSJMdZ9nTVLNPX4zYQ2j+KkBgAQjIYGfqXW41A0w
H2u+imGoWBCUfGpdhg1oCMxReF72XFkrkePKkpmlWyMYdVO3lbeGa9RY3xYHjKy0fVGBTx5WJ2Mj
n6jLN7nCH13BcjPsTpiqUkNl4LczHj5UZTmWvgk97HL/V9WtWzYgs8c0F2fKMzLkQr0hM+P/isuF
FIVI1HveM6jOzREM+Wpc06U4ZmE7fkqasZCa1iF+l11mlHj0dgUjmPF9qBbbJpiZb6msTLGg+TLR
L8uvMpwBT/vzaNXmaKy/H4o/KfSLdq2yHLxHthAhQLc6r/JgPedIvTys3I3hm90j8R7yMWm9rbx3
6fievzhvQRbTvGA5rrfYDhgj67olmQIBvHRlfxYhjooSSMp6PirUh7baFV/4nSm9L8PhmBaXpe8v
ikAyhu0KFEtg6jLm3B/CZ/5yPixaEO8OpDYuEhEGDp7t2xwRmiRoE6bwGNZZ0mZdVX6YvK4bSWoo
H3ibcWnuacBvXvXIUE+iTNTRQoIvdjqqCokvm75Hb9OPg0YcKuRhg/eM2M1t1WS6eQMa3a0AwNyl
H3s70aR6pBFQeEVXmMp0jHZo6tnJpMd/HrOjqJy8JoOa8OYeF9ID8UPXMDB+f9a/nayQkU4JUha7
5mikITjiXSu3P7tOyjzl/0SquFBpCT1Hq8lf5DWmIYcNUFh6Lthgqbf2N0E+fxAmXM3F066UISbi
4144FgpmiqX+Ds4BfdYdjwSk9d/zxU1omFqqurx1n3SAqGjOfFCzWS8xV41BR1JlfP3NOS4LoML1
p57IJdHMuEeYPBrDbMgnhn/Fl/9WqE7W/FQHb9Ugq0qiPYMigE2JpE5LruZxZojhH5KzK0JJRgOc
1JkYxsYBc9LQcTFDEuDr8pk8/boiI5WCZY90f+0Jr8er+pV5RMddDzWjTTHHmHuWyehuQ2+BTLg+
IXsLyFu/z6z9M8z69+x+o5n92GHGxmvK0onS7JuQ1kSlTizrWNstoVll5bTS3mGgdr6fHAGzTH4D
3WbYr+pr0ljI3CGNLyMvntTlpz1HIBdzIDngypMeSXEaah50YH9bhl5VvPncHyZ4CV+Ps+jRRf3x
veH3S4tLOpifiqzjNAvjlW0m+Rz+lYGJaFsRcBM8KInyCDo4z7ejfxmHmN84iTNhX3Q7d9Pk6nXH
qhwKXLGX7Y9YBkNncUAQzFnweyAINMwZYNqmA+JEyxt4O7Z3NkhKqBlCfHJD8Lvnx/1HtguGbctr
vXujxTDyahlHFEAX+SMjINrVhi3IMqXc2Z4JrYBM1TUPawnG+2RBVyEjwhVpqngxXM/rVbdgzcik
XZu3EbbG9SgkCBE2SKpHubSVloFKCTZ23i/HNizUkGQOQEewCTd2fZ+xXegWE9O6chXyjgjNrMHi
cFE6vazN27CUUvX+7p8llMstx9O8ZmWWw7T3DEF71YE2gDm6ITmBvLJc2x1PowVYOFl5ork7f1Jk
SyzFAgiVHx57oDd0U3HHkqItymb3ISEVdc2bW5sXdx1z3oF/0ayvATufEmobwzS6xiZ8g6qEH/S9
rqviJaW/tVRsZeaiz5YtcVdQRdJisEEYwDXTaoUPPyLXed4+KpcVFn+lzFwdRvwhXLsoEqoNznxF
BhFaN7vtfeyiKZnjtLa02NhE4l03qz4/FHqK++wPEzSe7zJvN4wx8UHgrNZFsaB3lD4rCEHV0llh
PpG+lPjfQud2Fjds+nQN1MhwqTjrAomMbWRJy3JRiT0Qp0VpfHuZEjcbJ8GdlluMFkK0rpSadpsj
cPYoqX4bgf7A3CNlBjfzNiA0OUcdNHEphava/InDjrAZFJVIk8vuXxC+KU5DOEY/xaqnFLBpg23D
JXdaW5O3xfENHjzbmWPzBuMufx59IQ/nRepyUbeg7fsgXRIPUMrXMfq5wvD3F1cnPDEllvvFDFay
tjM6e5hDWFhZydAFaLOtbloBWmvuJKMoaLayrJiXOr3GZNqxjo21rQ7DL3NsdBLYvdrL1RloToNH
OrbKdsKBCyyQgCvRKZPnTHcM85LptzTRhq0LvBvV8RVj0NsdsaRi7g5Wqv6dkTGeE5Rt1HkuV/aI
PbrXfztxHQHFjrpUi+stfV3EvsE4P75tDarOavjT4P7WUdadAoMpr5gsBKrrr/gCxfwSP68m+1Z8
de8GzswAw2S2OFvKRsbNt0ZQ9lIiymVYT6UtCq8qVzthF6lk0E8ZPdiq5aY7er2nhF40+JImYO0h
0DoTC/58WYCRoBU/UI0AQBtyrAV9LmrIHhi6zxEB2hbI7IY+vmTS6uYUONbKFIMKxnRdkvgM8VUH
2ROwwSbROA5oKegWVWRuWmOn5fnvWo8yI0LDFZih/l0eTKMqBnU2H8JycVG3zVMaJxLWpQ+D4sOs
xNTdpMTkSVOZ2CkSbaChFKFjFTaLJuCih+0iF6EXLXp4MqGHLSXdZq972bLF0zDyYd+7j+AIx+bY
PxsLt/m9DusHqXLQAbKGwRFRw5zf+wo0BBV1NAgfZobQjFie2K4/WFhrC+/qr6CBOIMvDcf4CZht
imZE//K8w/gqd5VZXgMO7u9Cn55y6yApmgCkpYV4PwAVWFzwkuv3ZMR+/QyZ1tYTI2MkLlCsS+dl
O0CZ9/WJnqWGF5h7D9VeZw+vAWPcmDhI9l1ZEYBDIfY76fCluHxWW60px0n96mguMTQobAXac5SV
2pKnCmsw8UZogMkc0Yp8MisJ7Ie3nxXpCo29FnbRPMJ+Rz33bgP0936hEf383gOjZIBi0Xf+SwNn
PItvp2NJPOWD+euvkltqUFOZaZJ40d2GeZztGdHC1m+P7JJOBhCTP7aW/JgDtrJSJtivKrdjpdMe
rDj7yRojWnfnVAsu/As0oVpgcvim1TcR3RNsarZhIALm1MOo+HAQghUjObU6LOSzoimUVi60hlrz
Ihhg3+uua5RGgrQBHa5/j1VixT/ll37ziUlzGQ7t6x4xyZaNC4+CZiI5yG24S0TAIIl9Ga5k1TSU
u4+Hef4NS08+r41id0fUqhPvf8PUx3Ihte/uE4sMCVC0haq2YnenJy8/LXdcQJhw2uOjUZrjef8u
abVHTS31DHHIRa2aoXxGyyMBe+2G4EZocDvnWPxTcq0oIwr1IIDoxW240prAKqRmVATLO+Wx4shL
4sIhPIgdB4Jc7Zr4u0SH+VEBod5P+facmd/klojZXvGtz4RaKY8g4DiTKehYlamWU3B1dxyU5H76
BlGcssD2p+7LjZ6qBBnCdqM1NJyWzjQpkk7B6lDFkUo9H2wW2HjCMtDNCNdOvqlxbP+EEE531drT
SnxnW2sGc9puF9+9LwOWVmkTKBq3ojaqimMMvzTAk5o9dmwbqfaalsYEX8m1UOrMBBgPt01N+zVO
HWiwrU89Jsjl8SYU/UQuMBYFSpmylTa1OTGtmK3WrhlI6u6+h53sHOh7cDkAMnIf2zvVKy7MY4xl
XJl+Ty6Up+CeXpgSoKvhpHBUMw3v0gS1nyON2nfSXBJzMwt7k8sD7SSaeZ2IhPdwWrliKnKKOg0z
fWYa3+MO6pQXoILGxFxFux6fyfOi9R36VsQd9OQFM+nn6zmCNLfvVMzjpXb8YToRr0stz1nINrvr
BfcJcG+mvjyyxaUHq35f6ZV/q3GrtwgNOKrwKuqzsukCHQTF9Ayi0Rlf1U6YWI9hSI8kJuOe4J8C
H6XRy/i+BgT5sjm9UZ83FxhwNtClwyCMk3L9H6kyWX997P+k+G9Peu3n7kxjOukbEfTjmhy0bkRP
7XcLDcR3DL+RPnYQYJR+QVWRZbZKYHtjrQYLCLiPwqktzhHZseEyegfLJEK9C+2/lxRQtRTY2kbT
7RJERBkMUX6boCX7xAG1EojteEaPfXeULQjN7I4sd4FG4HMGNdmnMS8StWE+P4JuOMLGe7oWmDiO
uDvFVV343sL4BuExOtUpoLj4uJm0BtGigH+Vpx6DUrBMPzYFXNCjWB730HCIntWuwC4mVxII8jCL
BHm0cgA9vmzF/etMmoV7csuP0ISxiOhfRwaQt1Us7Wmzrl3eW9sXeCQ7PAm3mMwdUNXVKBxECuEx
2X1LUD7PtRZZSRq/VjNE6qkOya03n2jtVIDuVp4X2c3eanmmszFyL4g/iAXRGgsumIBBw9qQkTQH
+sLDnMiDF9PNMX3m3Hh007PMP3q8fLem+YDCoZzsItGucuHV3O7MNohgMe7rJAitEX9YiZUWn18A
TCEr4Z34CscYoUGnj59XD06VN6YmNFFJqr1aWg/Q3iFOxVOx3ATUhga0D11aWR24VuHCjMH5Ko9q
/LmRVfcYV2eSVv3Yj3QtYUomUEE2bHlbyx7GLT0yD59Ma1UPGuLlb13eQ3PdScKhCfwlnv6RldOc
gggYpSjhr+Vi1mvnvux6YICuJVLuJMWHS45QEKQrBnQ8RH4wGCiUvUQuBZ7sp0oLWNjs33ANzMoo
9uhTQCtbHqwvs+500HAgCeNSihnD4gCd2ny471+iDLlwGxK9VQsTHbWu8ZxaE9hficcfKHZuqXfU
ufaDnfcT4xrZ4tXNBgEHXU7zKdFwVOcWeJ5P0IwrcXIOMr5V5LPLUbEdMEsUQJl1a+qnvQe3cZpG
YK8vzuBw5GvpTEJFe8ZDkkaj1S5tJ3um5elaCfSuQw/RepWtshGOnBXWIlTur+iuA0xkfDQAoEAv
PsaTsQ/9bYM4xzvcIK3xTh/mWtWDvd79YIX4g7IlWUKsWM7ceiie3mmbGkKSFbQtFv2kXgudcIKj
JMQPQQhWfRPiIHZqRbegLqAKMEfCOGEiLzLz8W1vtrH5SyJRhgWACUvJIq+AaOUOOzdX6pUUGI5F
oVXLKu81XfXXHes558bcq8fPoMOMtfku39JHwxDjdkzrEyIzqxkj8Nd+iOH5MDwOuMiPjrm1G42b
Z2ln6wyddDyHg3EN9wQVSsuIh2xT8NDe04j/iZD+dXBlExMWK2ACMpbn60wRt6efCeQKrBiZ2ocU
qr5yOqKSPl8oEoDli7wPLta5XQrEgxZ805dxp5YZO18BZTxoGuFgfgiuOFyudoLcv6pmtrM427d2
pKvv0px13btR1d4/FfXv8xyqfNmS8BHkzmBVmmZQrhnsWuaPDfD7QEtx+7aSZJpZ/cXryMS7lgVi
Bzxs9SjaeuOS+4YLFYpQpT8E204n2rMQIA8nMVuQu1MIzUROhxDRYo9Ee/IaiqCEcthK2J7SQRyr
MecAmcGw+ido10l6xe5d4fO+Pk6+iB9UzMxwfafTEqDHCvizhsHbvXmJAfyR/s3bAzGmScRuCg/e
GY5Gkj6R4vNcgGGCI/jXGQbY0bwD2aRiUlplMntZy8IQ00R4bMnqcIoImsXeTClfd5tg7Mgdimy9
czjQz7L6T1A0lB9wDlOeixTFJmSkG31kq30V5ionBWqZ73PmWKp1+yvXE0437y6KFje/vIecTHA2
H8dQp/opXvMPwdJgt1CiUHSKj8f6aZ/RvWKW74FJgQoA9fJGMhg/YFVX7apstbfhXl/zDCmBu4yZ
SQ5gVuERLKQ/4Zf8F5oLwREPokK9h4y6czwsG0fn/FLMeGP6elikAOhAx/F1HdWxn4XfNU4HYtgp
ivxffQrFmzNC96H8C2tgOjC1NveCxIINXlfNPQaTsf+A0VX1RSoQyqegaqIzOG5cNmciOODQAmD8
dKAa9cTknDxwnloZ7ozLr3yTUg6tHCyJ5ZTvWQixlo9m2o9hWKFGwqqusALvCsv1INYAzD0hjJuX
zsj7WKsPut4sjQEXP1SBRbvGKkcU46x8m+FFvHneBOf2vE+R8h/PrSlOXUVVkjFvb1NoylIDp5KZ
4R8dP6RnHvooYClR9nfyi0OYVDNmlGnjGICq+eZpdEcvHJ9YiIUX9yKLILX/8qrIb5zysD1s3fKC
HWx/qQ1W4Qh0Gz9Q8sZ2+L+kagrqnkGIbXs+JKOjxQgY+z0DaBK8qdV9m92crtJc7exdlthgdHHa
3ruaprJcD4toV7Ab4CWDhGCo3o9+xAM3PWDzq+0DYQEvAWxikhl4x50c3MIL9ymYCwhaNinWHQJp
dgcIzoG9E1kmka0F7l3tTYlLBaDfCDmkmrWzWoeK36SQFkJUE12jdGQH6wEvTnpYZ/Ost75cM0bH
4MK7C0KPkAvOrlG3gwd3ZE8xvfz9UTuWKC09s+3era9+vhA6BwSFhaw5sNta5ZwSROOFLkulvrbX
NvW+9dWvDUw8dIE58fZwuMtqH8Deva6yUewxqXpHuZ7LMXpGYYku4ZRzy2LD0CYsd14UhPWS3RyD
G8NNJtYDq3YzGq3d8c7mJBtI3wRkn2fChutP8C5G+6NYLHc+s44IqTjD61PTNMAtk5YHCXJBIw9y
1QE6wo7irsxRv33tbdY6bL5ooj4VtofvZTpsNMV/E5mu8kyaeZbKgFFWPuWZRsBblgT5s9lq7lqG
Xf9qbZU2W6zZngCQ1UN9NZUHg1hxjdozZOQVPdWDQJtheYoQMNR50i4qehSXkY6gCVfmpd2jfxYv
cE9eNQZMIwMdiEek1LGErY1VoHCW17ljwkqZwxg0agtUHdv7L6a63ZFspudxN/f2RjK13Z8uJJz/
2yqI6dzLhdL3iimQi3JS5lQIRphQgtU4A8M8zEmi+YrYi+TYRYw5NzUeo4SmcQ9J48MuJWkXtLTu
y+Y9cGjXVHxWUglURpilXi3C3JUb5JH0vy/NHfhs/5TQpAWJ1ts94dVaJNvwoE09+MVjOldnsoi2
HOWjQKeUZlbFx5hoQu0Mk7BgezBvRrhpgJBFJ5rcJzj615HSLjBlSYU8vst2jp/jNBsOpVKAlxR1
YbGewWxmHwVmVkCRpoKKNTgNKwt7yF2YDsliD4yRFRlW7TlRbNzFj33L5B/gj5xaxVe8SSF6xkh/
8mPhnywmYRoNOBpc9wzwPhMFGDzaRx3gIz2M+8z/t4O2h+rBBau9ed29dJfCLUXXweNvLtxK4+7w
lyiqtoqcqcRk9JfViT9BgXNksLV3sJD+57FzZnWfI+uh80P16h2a9wlpHNLEKK4OTRpPb+vNZPEw
88QrSkN3Y7yr+53lciTpBfrydId/Gz5FAPumABzR9c+s6dLgzkn+hsTh9ArC4sixLiCGn+FvK+Je
x5LDXX1+7elZqnnMoNBvDRWj/J5CL7dQcgTL/wiR3RCkaYv4LIQ7MOjBN4D1y7S21QUaLSBeCio4
sfLRG19TbOs04ficb5n4H0i5/d4Fg6Wi1huUrRt21449dweVSSrYgc6Zye9TLhaTyjQcZ++SP4Eg
sYhIScA85w2MGlcjd4+8WgGBsJZmYEEa3MRlYIRSWIcpJelLptJcEytImaoisGiHxBLVZvcHSUey
qADoh7Zj77fCtsZXUs/Vbnj9fghkKq/DwzBJXTd+UkLNi7pGi5xs+aUUhC52DOHSY6jRJBClM7Cr
cDZerdpV2O55Ia7echtxeJxQR6DZoyMYjPU2x4RU+qg+IiscNdxNLNEzeqG0gJuL8+1XBIZxwXKU
lnwL/OCQY+N8sYfPF9FlZgPhJ7Q7600d+XBVg5/1yT2kiRH6n7IGtwqYlJeT4HwGO+u41cd+MgWv
HkZa9EsjRhdQQfssq7KUW1QU1dh9EgiTl/51QRSMdn8YLRvepuzyrJTT2xPzCecFfmsCFYusBBMZ
eXDt+uTgLS5KvDogF/e4jDBp6TeyhgBWt20Tc6VQzXhUXQdFE1RTfJKAmdpOJqm+7P37xLVclOG+
HfCc7CR9Uzkc/yr3/yYdin3GtX5Juae9nnvKi8MJf6DIfDd8GZ4bPNZCHkxFtzEQVGHMTE4syPSb
GDb2zDF96CIqRB5WL8QejsqRpUDw6OwcUoKuk0GRlRz8qG6ek1oaM18UB+IiOndNFBHY7hfBGPDo
0FbcfzzKfarrpVR1on1rrouMht79rezWdb2Ae8FhWf3BNVIaVGBi7WFgvSVhChUp/S+AVWRpM3CY
CrhmMlQb82TqlbZ4NFCGShL+rkHHxOd2cZhaPrbT7mR0lM3lRfKVxRpn+CiJBAm6wdAHZoxkmT5K
iiV4TI1gQ9c00NST/+e5++MbRY5BnLc0fqRZjtU12sGmQWAo1eY4DAPyMWvPrX23e8yA3ofFuh7n
7Y1lALTvHVj6nPzy8LDiRBUdpnRz4XR6xBZRxkdWS2AU06yl8BCOo1Lj3CNncOqxcMg+vtDZw0gV
dZdTifrryNYeHxLIo2QeTIXV/Sd0kIYO76ror//cVar/UGWN4Hcddr8Kbj1TqbbVMxdplu5FGPmT
AjvBYc/g5aOLAnjliaz2UIN5PYw9piBJVN0Ciy2HbVywH+LxZe71L1wmcEcG5b8ioziH4AbPsozQ
fQFRB+tW31BsjdZgeyaRfkCHr07SE3rdG+89EkKTrLTBa7RpN0Nx1MY1UUd7SnlMsKVu0Zy18OCo
nyb9d0+8Fd/Hu2DtIFZ5HqxmVQcVyfufIuVT2spdI4uOco2v2ir9t+1gAx1oHmxOPMY8OAqtaRyl
YQtmYKpu9TdfBmuPH6J6agXwQ8sfOTrzddMYUWTEOM6a1WbjiYYFFl2mmShnXEhpnsA+QxBcYgEP
OJrYnIxd2EDNixzesiDJr5E1OwT1P4Sppp1J1XvzQm0JdA4Fc2Wqj18zP/M6keTTXy8drk9HCcPm
QqYuce4Ef2k3jqDeEDoBnMv16Y1dy5h9Su+tEYAoJN1E7Mlhu+R2kwexdnbbQg40zIv+H5xwEBGQ
ES+lBFE++cgngdC1p+T/brzD4gcdYrszhNN8AtHM86FArZPOXU7+ROFpIbxe2CUZR7Dgji3nYcOX
yzCKp1Y1pkaGI/OTOt8DjiDGurl1GBjZfCKky9wkSqOzXL0dZXibOJRLltKZWpREBHH7ZXEHazUR
WVoYdYzhUMNyrl0AkNKalBc+yCkqo03J9JU1gFZZthcvsseudxm9x3CXoRU3Mw8nh/ri8YyZGDIX
iapbqU6/Yo/gFu1c0wzqqATHM5/OQjs1n50Ej3136rFjh1J7bcDXUAB/g95/6TU2/ypefbz9JPIG
usmIjJ00AeG85+rljDq3xnFSCPsjZGjk2r5dSaCoDOzvSgdcSETA9ULA4t3ucqH9Nm+BEwHvkVr4
FqiRvZsUSph69Cs6HVxj6A2evYH22r/Iu+JvlYg/wlfZZ9y1R4+ckS0A+++pidyUYGTzV0ickJuO
N8gPY2zKKVgCNY0nKxYUQA4G9Fc0jChCsxHRJTJZd7D9NuPpZOo6sSC9p4fdu9eC/kBck2tCb08g
zElw5alQLDCshNMgXKjmlU6zU7hah4WORXj04Onm3Mmvbfs4rA7UZLFqQAtw2XvXx5OJHYVXMaG7
Gwrst+75I4+D8uSC3ppkngWGvAu2tpskG5f2TJQ7X9JaDGnq8pL8DEiw9UKzF48jblkaZObTWD49
K3XfIoydbkBqhhSkRwCzXnCwjxjhq3Y6HQvWakfr7TOaR8gF/FOI0YCEp+3YLRYV7E61chR0aFAF
unO6IP17suc+DhIYAYleJ0H1vPR/ZOvUA/htR1+gzK0ArBOE8XWjp+mksIWD7o/xmQieziPoKd7E
bgMSuR7AoP33iF8auIvMeetvUWVKD1BDn3D60YLu9fYHPhwuObub4COm3AEGThMj3gneg8XD2Y3h
J3exF4y6nMojN5e0wDtu73KqlsA/9k1Ip9t8Dd1QMd5ZSQU/OlTm2NhJ42/2OVu9W9jvvJeWtv26
7PoKt3LzvElHUiX7tBm4nwdHHzYH15LoubYLT2UjrBCY1PCsd+rmQ2dLGYnGI/lIdIVzgVYj+MVS
//O08CD7xTIGzEiu5veZ6wzdmQvEGCwfi0bHqStFAVCb0uUrrworioNOVpV1jYb/CUdOmovjOxPJ
NtFvU3KVFzKCf1LOpqkeXQCdwe/t5971g3T6Za7Mxj8adnkbNO5QUPXvvGL3cuGrbWazVghWiEDW
9P5bPY+TJ0kKU9T+sG9uKXa372GERNkOZiEWS5wtKG60KusuDG4AZw16Q8XH+U/ahrhzW/8JBUiR
2szgcyUL3PbVvdpWVe4S0LRuX0rXhpXrwIPlf7Xgr6GfkU43S49cJitawce89QUrXg8pNTU80nN/
XVzzFKWSpJh+7VAsocdLqRtwZtJLdXDi9zpxC0mP0L1XQSe4xOiuyEVCqfLOfjYS/lF/aQXbk7q2
Aw6CxEtBhCxcg72gDd5xQImGFWR5UcAz+erScAjAYv5kkbyziOliBYAC0DQ2VPBnqPYVlacVD7MJ
s7CThTAygXbzlnydJOjj3Zw44omBA3eYWVPbaP6OzFgAYkSv6xvzFIozQXgWDH16i1QHPc/QkUbE
bcM2QdbIyCGNTCqvJYBmFjC7oMMGt0KJEub9CprVnSdCAJ1HmUNxcy6UsUY1BhtbCnLiKODdjJ3N
hdxccdWxdb8P1gHPsIymUDHvYGN/y66kLcMEj4QRzB59UUV5XZ/PW2zy3xgLwxJukaxrkCsWqYmz
gctuI5e48t2MGbh3l4e7ljSwxes65y0kwZxT3cTo7Wp3ZLiKBPhcwFqMpOD3839uYNStXkYrZI7N
c6NZtiTSuBQ168cZUSjG172fkrBKuMnYGz8iISRoafBifnMfR6V2k2yYklsuv5gORlEL53SthwO8
ZLd16a9MH+ql46lhumTVYp1bH1VPYuwdv/9bs95dpCwNdJLlYL5D0UEVJ6c1ds5Pp2mi2PF/NAdD
9afqdUizfOmjT6kqpzaC+/22nns6XI2bh1a98q00iByZi7J2FR4K0RgdTH4EOcz9gOhPFfcmPLjV
gWh/zuuulTm8zvHbwIS1Hdl/n11I2CHqv4txzAu9lEsebWRZSO4TxbGm35y3LZ182IEcGC81Pmwt
p9XzyfJeXzDpdkED0W32ZsF8Hk16xmwTlmKsYJ9o1iu6tjKPzPl28TjH3bTDU0ngTvCSRAVgwKq4
kjq6fVtRy6G72SX12NuqPp8oaP2a0/bOu2bGCDEj4fb45XQpJWoItf4eeeZyWu41vzkE/b3TyAql
F7r02MxUZ1/wthGTCQKJSWufGVTrFTbViLq2nOymR0NL5qV7lWK4nV8Sr3rkSN4Xb+uHjjiDITpX
FYlFH6n7Q28BkMj6n3W+yvVo4EtfuXS70aO0VCat90EvECGe2PZjIfYmamOrBj0PxFWFLzmdMSwt
Fj6yHtrfy4g4Vj5ZzIVtvV7nRpy81SWUBXI6XXazZVbyZQsCzuHjM0d7NyNFiCCxTmlMHagb+jZV
kKWa8lUOlrHacBAjZlVPDCI99LRfQHj/gtuBGEv9z5Xnnl78jpwD8kbd19MXdaQ6rjqyRrvMF01i
XFzgPsMNaJ6iw4UY7RYbzBTjGgIi5s4EV5JFWb50M5/3frfXef/80b9gsfhYTtbz0teRH49eOyoN
ghFDmp+Wa1RalVNznzu05pnphLvpKr+ANjx+CvN0Egu4nTKfjTKrZkn18AZebPIYiauIOL4wkSku
MoULMcwbqgKBeGYFQ45mdBs6xxGc4T9kTAw0oEntzJx/87G3qXvtiuG9pLG/OW1CHlMM/L8FQ5ZM
1F2CLZk0dRwq9A5KX76rnZPcCm08bh0wLj/AVKoiKsSEh6W4Bv8jcJ3DYjx5RqQhtFQHWMMkSzGl
vgovbpHgyKqMyrJ1jrDnBfkMtcsZdVLsz/ggxFywpl7KHS/A2uT3uEm7eJUfhFV+1t8H3LqQH3c1
ePd5ucmn5PKpsvV80O/Z+2QUd0umyjhTkjfh6cGh8odl/ZpnV5xv++oYqEn//waaRBSmCOIcviwD
jz/Dqwbv4xlF4rxcee6CqcppXsi5s9BG4PIOGIBOBAUa39olq9/CdQ2LopK0FToJI9OoWOHq5dUS
u1AkZr7SBDUONeqxqDqRtEiV/hJBVwUvMrXPFAogoAZ0j9N1ulEO/vubPDEKCChWTPMJCLw9XDOs
dBGrcpQ0KfvZIZ2/qNkyiI01rO8+aEhiVm4O/i8wdGmqjrPMvlIct/4xa0gbcFxMyxKQjDGj2bur
5nq32rT/Z1b6si+54x/J7TICnJymE27f/rYnABYJnkHXFKkB0xlBOy3gTTjG9/p2egyP7tHXICUq
CRj8Fb8i5B6IPZiVcYuJtKQt0WjxI/1NQBkaTEwZQmJxiXW5/yqywbMTS4Ya93qxbz//buoh/VT8
WDiJ0r0m83bfyS/aWDqvmAeACokYmxpVEYLBcY82/kKylcr4PjPJ+o7njmnr7OSLlq/FRE+TIODC
aQb+VkdgjVGYwVH+8clpf5p9Wcw0j/h9iNEIk5cL3saHet7yC1uspXOyEqyKTyGDEtC+rLKnolet
hMNjE6HpAN2G2W1PvOoDE7yZtcD45Wyy7J4uj7i1tY4UO4ZernLpRBEB/HtjFpxboslC3aV9Z1tB
p5+ao67P83Z5UK2965RfcuRFcq5phJ1HgJ3/cUFFbpcZFqUfmCG5QyPVkyMgr5hq+gz4qY+7hcmU
94TiCSx1al/1IwFOu7dwBDzEOPCsixndEONd7g3//qEgKibAyHEH5wW0uQuQ8HIETQm8BlxCvHzp
TM8hP36gp8El9yaXSr+2sQb9n8Y7PPaC5lx0tVKQmMsQZ/qrf7COHhbZlf5NmrrTuqHd031nk5Eo
+tmdj3bmP0PSAINfWkndmTl4E/p7+CEaniluJnlAc00Xh/T7ovYmUWOBjXy398zSfeT3SvJ5fU8S
FLur9v6/6v5JCfRDAlr6era8LSTdgIZARyiZrMEEcuZZlVV+WdZSzjwVvWmK8/EKUKr2WlLG0Gis
0UcCzVW7pwdfp60SMXtdY3+7GxBpLjptx7wUSgodmmzByg42I0V54bFcqAHjurc1LDZg0ge8fNTy
YZvsrShrgqSQjlzfXjcuz5nue+WWJc8VFiiHYoxkjHa7omRFhBbcUHhQeGSkZ0u0/AA/JInAHpzx
Oy7ralIkVDL4ZPUD/MGnRGH49aQxTF6owGfZl0a8pybZ4r2/Cjrp6RWL3SbUWOp8gEcFNYV+Hk+5
JsbNFc6LL8dytHohdw41nssoALkfWU7/mFVbrTJSwDFswAn9tiSaNibkJrfhBIUP3JW9gr75mOEB
AGAf64wwlIBJG/sOKDaFCOY2u9BlHqIy0Orl52PGproi71uflV5QJHAbSQ0UR1lUdOBEddJNvEe3
8XRjwXfCdfUWbHZCXhqpvYKnQC/NmY4wNlURVRJvXdl9GHCOz7GjOTFJzHPvTPgfJYQgab8rKHkN
+3bSrhWZtxszf9lUrrVJ7M6SgN93X7VYLERUg1/4nv8tScqrBzdovj+F0rKT4WBQu2VDFGwkBQvt
7lwrX0pFo1I3w7T2pzNA1/UUlo5CWuP9kq2jO53wd/3Jg2E7sVPlPwMoINUcV+clMT9InXu/aEFE
I7V/lHya41WG6B7hODg7G+XCu00cm3Dyh/bg/MQtipV0dYNuylArVIcNAeBDBV1E7GwwWcAEwbr6
xzov97qL4HupZI+LDGKmYLP9PnWlHQJv3G1Q597I6co67+NwEhlr7vZl4o8KHykFKr3NoymdIQ8T
daHl73u/V1Xzn2fKsMVDpXrLCyMK4XClSqpFcSeauXVwfOSHK8XVSxHk/BeNpefDXzeaH4A8aaA0
7wcWAyquP+0zwIlhb2BQShFzGAKyHuYPCo+5BEIlf7QD+1gMq/XlZwJdDGO0VQqNJP+YU6PsgnfK
/n2htYtCECHGL0RtYKDREw3K0LV7R0U4kg9aDVrEhN1SZhlPXq3VV/qBpCptoRWcGYPJX0yIzH0R
heKP0Q/E71kKriSt7WWTyda/ayiM8+O7Wo3H84erUhvPQ1KnMK1nW3HMKtpPpGEf9wl4OKjGhddi
pgz3LDXEnAG8qwZl61rnP1GAY8kbmVmp5/5qRa3yclHJYtJIOju0c5JYR9olDGPt9NnaOgDyJlKm
bO2UrF3ubbfAVOM4Uc7vqTmGZvQJj3LoVfNlqGpVJ+cYa6x99jeGcx5RBijPXmmYpZD9OvzkvH2+
B8ijoM8awnHHjrybWsb7fs4xcbLimR3oCtJz00MDj04HK0o58Hrz4q6bFa9Odw47AGuJQNnFt6fm
6/tcSKAWCw8Lj5uuCcj1mnGAUs6G48RNu4vTv8g72ODYhe/QkrpLJ3Qfa2oyIm7b7q+Mahy3XQoZ
P6HXBjEC8IDSNB48j2GfucXhnDI+axtexlD15aBQ6nHSSZiqVPKaXnRN431rBkfJe6b/9Ms1wStQ
rO5u9eSqDDzx3Mw0mSXmQUEMzaQC9b9hJckCtLwGtdrkhtarXGb03fg676u0yISTSxNmDvT5jzbL
EFvnK9YuEHoeU6rMBW3CYdKFTlf0HiASImGB8XJXuxEltPZbWHtFUMv7nXRDvlKNhrfKCI9FyK52
WGSFc9F5/WIOAsYQaNyKYGCow+09jzNrnfXa4U17lZsaNsaQFwaqZ+C7n7CFf2HQ/gy0knKQD2Ud
M3XoGp02WI0mDvoz5FY8jq7aGr4u5VsW3sbvhNI/YHp5/nW/axugL1dtJPG9HPe9Gg71za6rThnk
kexnC+emHfoP+RH5bbeY9HNWczgRtGBh3B9I3E2NhU43scCifflEpvJl2e8vnHMem1Ov4f1t48ok
Zf8hdfXX1RP/cY06xa0woaZTBCteXcjQ7LodhPAEC/PNAIMkko2QX6uI+CCWDEtzRX5QoCevoV9D
7O/c+H1WfJfC1DjDblfOnY5UXbbxlMPwg8iPO3cKKuN+uB8+QfcJzj71n0kCjSuibNXOZ7FWh/GU
LVZ4b/8mha86HgAPNRD9rckvHFVWR3Rfwq1iTOLeDt3Qfcb/boCOwdB0swhBoBofakT/tTdwC0a2
kxy5DuQ7z1kdSIAOxntVI1VW0Q0KwbZE+PYpC3pbUlri+7qUW+HcBZiw6hwHhKrTw1HJ++0xBhGV
poQGRAn9uDaZFA51wnPI3Rf35pCVpD3A+d5pXgtDVulcphoGK0PfGsZ/5GCzJLRQhodzjMB9c95L
VkX3r+DT4Ik74YcMBLEgaj/vq+/tV+jhPch6Zc8tq08GwaPklmcm0iRZJiLRXs0HbXGiVLMvK72b
d5gQLFU4VwGDvkeqSzyIxQidGsSMZeOQBxnVT8klLvlVMnugXA+16lyzNPC9wB8oaubPG/6EfIVF
xXzQuZBjoqw2LOhl+OZpSpM3CeXBmRR3YHC2++xQQdmzaIjDTThcPU4nYMOyr90eZsEvvWheZ0e6
ROYutFK/fdBv8H/mD+RY/WpBEXeED60zHHaMbyOgRTSUr0ibA8MbwGhFW46cScZsSDSIG0Fmt+rf
iCjXTpMuXXfvwmyZoGySFHydPOx0zYd5VgWHd5O/XwATKl1C1TVOscLNk9N8a3LWQ6xh3LOaybHf
/ZDp0yS/ZVtMSf8B/xnOir4PgQQE90snLr4SaJEhrqF6Es7TFQaMAnMF5QVe5Cxd0gMPbf1V6KvR
PeCK6g6es/vwj4afVXOJIC1npRfP3LzBh0oIZLCnQnQnhu+RkWadPz+AatyDuzztqmYxGl3IrA3y
vx5ZlPyCPSCGbxvR65xmJ72kz9QI5dYYcgghkKCX4fKh5jAQg/tUJ9VuhajI8vlYn61UbNtCwFXT
B3B8cTr5N3/4qN5h8ZqNhsWITHQsXfVfctwlEDmWpyePn/TppnSY5ejVzajv24Md0xFOJePKw8tC
Fj+ma0zFm+aPfAeOsEchdsFudJVpW30IfXjPAxbAV6vK68Rpd/WDwW3bTmkD7TdKF3r0YE64B7iu
bTeQ5Fqygb8QlVbEBq62bKQQwE6siBkvgrngSzHl3ulTuWi9PaIHdR06+/cnI6TTDMvhNWQIwDTj
UNb7HSn3T1fRRif2XKdEg4J9moyGufTb+fRHYZ2QNkrW+NcU6ZVm0k8LfpeJv4ldvt+Gf1Yc6EMA
nXHOUgSnscU+vK0LUAl4rJAEMUEmbcTKdeMjDTCgU55oqKPnqFjCH3DJB2cNbC8FuwueocJ6sguo
B/O+oYaOEMMFiNEIbTD51TfgA1OKm7Gqx2BaxeP2OAyzBObWC0xd7iu/hXMajTkMQZPBHhxTYlYF
f2JvuntTXJXOkIsK7YwlPrqxXrooMRbIzKwUCu7CNacijJA8KFy665tIh/THXAIqOhpZylhzYWTl
jrUhINbZ5CrYvvHEdXCoEbmdqhYx2kA/FOF74bJxjQY/xphMf/GKxanWTWuod6TKUKPCH4xoQtpv
0vJH7UuLQUy5CU3HF7TqwrafulgoMNrjbLhnHgdi95P+csZIBT7pLTsQ1+0qZ60MJdhR8yhknomE
vnlpa4O8OdK4uopWaqTi90OdBEvv2Yb/HftUGfZOOmT2H2xorpEA3+ab3wlUt6zGEUFjc8kmjyeM
9QVtKC8ZsWPf3ZNAtC1HhIR5a4be4zZ2zkwSpBHpURvQNOC1bYKCR9t2cZA6gpxpdjtWqsDiVAcr
lgCgeEiJZOvY1gzWAeRXXcI8upr1ApfUrBbchOP1AMav6xMmwHYU+ZlPQDC5qSMWKe99K7CPLn+k
5QekNNgIiKMxvJ8juCsLHda9pg2LD0K1aglntPEec/jYMYFrkZgRAG6C59oCFFlSwzCwa9cWuMx2
0L6ORs20aNvAYEUbTWW2DbaElEaN8vTtt/5kjcoMCOF2p3QDIwdsrEF1s5DylrO22xlZIDvwpYi4
99Loi8oQZLS0YO9vVGFCDjQyEsnJ1Tj5KZYPN3QXGckSkQd7L2dibWsYcntS9oHKP4oCaMp5w+Ya
hVGEqQy4qkLULkNdFS2bVdW11GxyyiPA6eSz49iXntxYZwUjZz+wlwDrRlxqgVYaUJX3D1VxtmvN
84H1mnRR0iWh0za2hbJBj68N3/dEicTGMmAXsuCUB7AzYf2/i3o+VoqrVWQ1fnmRvap0iFIdsU+V
yGEivtWxEfKQ5GeYYafDDbxt1GAlVHpbUQIkf74HHpNUsu7NrcIu955nSb7ct34QOll6IBEUhyFR
U1JWwx88kHUdtYnJT1kRNEGwjk0QfZzMe+zvmEatgxsqMuYgCcQ1BLSIkFGVSsP1n4jo2qBL2xBr
iBYWE+ayhzP7TPlp9gtXswgEJN1HUp06YlejgNRScO0O3NTDdz2Hf6V5kDnxv8nTH8yJ9hVoTsLj
J8QshLTIdPtiz5pj4lCwDsKCMmNut0Kb3pT/HjgUAf1olzrLt2F/XZ/HHGnLDen8T6ZJvmuKUMU6
7Davaw7KsEAUAdFymoXldww12daxlqYT8E52kWYwplsbWqVUBV7UznVTHNsK6RJIsbDsLQye6GFt
HBx56UOXu/0FfIj11OQFQJipTyDeBo+KV1kejyIONv4bwpC0lk+TWnQBHGJqu4yulN+A16C9aBEA
Ecfm9RJrtUjHZAnTxM+nkysB4qhG7WnEPh+MN1xeW2j/biewp0sGtYNcS57SDFd8slNOnY+g3jI2
CwTP3mG9A2xLTBe/LInmOPs0KdyZBFFD5QiaPTGl8Sbux9en9FohIewQTmC1CJgzkFzozqnetgam
4UR3fM2sOtWNwgyUWQwD3kpAnhsvbVbDEqmop758w4yAUvuOGHqgcdI7+uT5tNR2DRoZB3GCBWOK
y17BDhIqvoOv7IE76Fvxz6i8gUqbF0ISii/o32yp430G+nNor5oWWq9zymDlf2UZWM4/eX2A8+XM
HYAp0bfh6WPObADCpHbNwxKD72NVulj+CGW1Z1Iatkdi9rNpddAOwrDrvXV9MARt/XRCY6/kYPkg
68O6KHZPgU5tLgu1W2ZkuhyT/kb73y7fcuKjSYgqy8oK9+VBxWeNK7+ZE8m5lQqZ9u2M20b3ys/8
MX9J/3y/mIfZ2KgQSXcXvSYMmyk5qguQZLCC+ZMSYV+zY0C6IbMtADN/c+kMYtV0ZLotS8nEKjD3
NUrW+nZNQ5QjGxx6nbtp7ljvwkTXv4d1GpKXuiS0UsvjBhmcIrGNN/aLAvXO6mVSYpg7XF6fPlea
+1WS07SBnOYpgwpzwPWeaF0Z3+brB26Tc37i+2X7A3OUiwnp2pvGzRWffl/PzJexxPaZvQtho67R
VUvfNsol+d86ZuxWoErB6eKA1IWOnIVlTZNzz7sSiTPvExVR5pajhtptrh4oUoDfTveekwc9vQsU
4xPckuPhoQ+SvRA0r65RFk+fgXGeDlh4oTP8hzOKDWqFCNkRnqoX93hDF50VX35TxQn558VoYQ5q
KkPW1NIMuMIhxnveUS6jJvbPEg+eX2G1y+fK1mcSaeSWSfPI/LjIlFeOlFaiLORk12vL+tNlFM+p
zHbkkE7mbaPB3eH/TELgmfMrdJnOATlZYCowByFATmBZfaktyKz+qi87GebGDHGobJFEkO59TnC8
Ce52DaBKcC0EZCE/IlXaqVk8N7LaOafV2xfgmWq6js0KJhY2527409f0iaqaYJo3vMQt5uIWcFiF
4r77uUzB0/ozHKboAley6lYLmzeUcg6Wpc0GZkfl1JtHs2w2tMMa0JdGtxcqVWIgbKD4pCSOPzAW
OfbgVhgIC/N0roLukcv3Y/kRi/MxzivkfGyqpYJoXEcp9VFj6mdPc4IXdIBMrrc2oyfJTJWJtKGZ
OHaT8p7RFtZDwSvnvPqfEbvMMcplMmCz4dl+fyBHblW4ZM1lPCgst4WDEh/uTanAlz4p+XFFMNnT
QB331YS25g8cZyGFwCOfcMtYUsGkDsr8b7wrTYDB4xblMw+VJb5NJhPMQsNKr/dosxdbjWA/Y7KS
1Y10IAu19On8djN11ioB+N478SAOcCsEiheg0l5aMVi0krvKhxZ3x4h6b9pj41HyXvNG8qUGfWpi
jGqC/vbehHXLKvjGpqaFoVPey7aN1hGMNxAVjeVYxBnGusa7QLOcSbTE6/oVjDVt1Kwr14ChoGLL
Y6rkJf9blcEir+Fa+m15JpT58UAchotDol+ftktH3JqVg8qjsvI0w4SM5gA7wfmTXC+nvLuzEU1N
Ad/iLHW0MU92I425MyqVQ12ONuWw5X98fAiCSr+KIJz7/KjGMUrsKVKDxyekQfvWa212ZXMBq3YL
u2fiR0MCnloo2ldkWDxIw/mUyfiow/XtJm+wN8SklzlRFGwIdJK7hhJbglfQ2HGB4/ZZ48HkcLHF
IXhNkWBfaLLORZGH/y8nmmpJaO/okGXx5Cw41lCfyWl56ZB/mhgzRnRe40w+eY6Jjf5LMjknrU6n
R7G6Ia39XyC0VX9aIZ28UUYcB2v1i1E3rMSxtBs7krEy5xPp/xuunjPeIWyPgYlmvK0eSUCaMroZ
EVyC+QEjmmPz1hkzcrEnXdRxTi3oeeBlSE8XlfCuRdyOw3NqqiQQ49b8s3jyHWDnZ47vwGtNH3Qb
3RGhivE5GCWEoXNQ3p3Q7wrtgaL3kfjUx5UsgiqAWvJSjQaql0zmOvAinYuI+ONuGPuOPH06Y6h+
65hqUu3fQbKJX/Zc0cTtNVux5v+vR9DOk13qlbU4omMAT3WIQWV1h1RYhRrpIIdy1H9mhGMHmonR
OWe1HzrTA6/b+nsIlO2A+zTK3mJiFuOILRJ8O9VCnDzIiMUfMLyyw1990P32SnaCS0vMy0hAUTo6
ZuCp+F/f0AHjTX8r26AObLmLgv/F+aKDjU748ZkaGLGajnusCPKomS3rVNZaBTjxtvchsIGK4AMo
o5VAEXhplQAp8vQ4UIvAzXlJSZ5ntlytUHck4BCMZYYMeC2elIq49oBS5BV9hNC7HDJ0nrulpe44
zaCKudb7+Zlnwc3gT4IeYfTNKBvcnD2/KrlQuBGNaGpfLqsWdeRZKylQPEAtLoPIMCu9psZD9ycM
2oBhs5rHRkidVimdcDUgqyGT3WS0olIbOCaCQB9BAU+KCBV4G0jdIuVs3zffw5pgD3xHu/C7xadu
px4+oFe+A4o1ipGN3wqSo5HnTWaRrifejYBFLLIAaJbL6hlQz/MvLq39R7uPOaifTkxaMVwWEK+c
vmFHAlyBLHwAOetPXS7oNgbC2R+FmGhQFPwfxpYS2JctJWfQ96+wrqFpbdqKStb26deRcGHMNbyN
VkT/4/U2gOee///HkIbnPZv66wvSr6MLib+0QsWZbVuKYbKcaEUGkLEBKLRj9YLuxq7yWl3rxtWO
gIuPUGaVcckpUubao6c/jK0ms+CdOVsPF/3xSbu/yzkZEwJV4M6GsKVySEbl3aFlxIzNF5XAM/PL
8OD1l7OvyTEA0HgwAjvTIcH5MZmuWISSn+R/36O0mgflNbSTbmhPdm7w0H5CI2+SpbRvxr2txE28
daTkFoZfwVofpMsXOeTrGE9xXF/mZqcUSuZk+Dx5MFcANO6udBwscqNdQh8FZDnhabP4lTU6h3Z7
mz+MiCXXAWKZSunAJnNFr0GYnz0au9hEWA1Y6ilkI7vgYCwLkRtqAwcVUVprmAjH7R2EY2YY/qxN
BPmS2JjF4uI72LOiM//UM6mkMCwLN9Bt7hWbJ4l8a3hyiQTiwJ3PonC0BatPy9487uovZW1OGIj3
ITY1rIvD5XwJUqT7+L5bDHkDUT82CEUd435nx3zQswYeATy41lCW7Xh1EhIcjG2h4vGDmMPpy4Uv
o/eF6OlnU8Tx+4hdqzuwYWty0tyw8aMPEPzicCo1hRREBLXfQJ9GLLdbCvNYMZlYlAn2Kvq1Y4f1
IUS2XEmlQ7gEh9zsaBhfAmJBiE32KCmAcr8KxCDe9AnjyFnJ3X2a8zNFdQ7Ubmq8XMeXCuOGo6ze
4/JstqqVuf+cepNgiivtzjn4XUQS7+4l0gTA3PnfhTOKPY8MhJ7KmnCojMKfNU90hQvIPJ/YwmS6
YnJYJp5rViIjbwbKceYQBk7o7JQGllV1H2oufTpfckcPwLHQxGca8qnOlcBE8gnkq1ii2Jd9d/9s
nMEoweFPvlrDofICDA/WAlMDcUqb0QFkiXK+WSlxrzCf+otCH3cf2i7bi9eJMkft8AXSprik2nHD
c6WChiXQsBPNdViJdE4EV61uoxG9uN1vjOUVOn+XllPZYt9bOgzccJTUx/DjkTPGq/YgwxMJSBJK
YOFMozX5s0ZU36UuvAM5SKmS62gimhLVB9EDxIMxPR50Gr2841SToUkdOGgO4AHjFe6zvwWmbrM7
p8HFsCJxt+8no6WUmw9GhouP77nOWcZTMkHQXOm//lMARlF9SJv/bMzNjXZa+rl5qqvlKlEs0aYQ
ImRJw85aANHURHcOZPnDvxK/q45NV2kF83KEx8i8RDYU5XYE3nEmGR17G1FHqDieUZN5806IExKF
njhmghKwc26SLqvwdEqMcO3l6qsy8duLX6Z0ks5pKderQXE10arYRoeSvB+3NtpzeBvX9q59WNHe
z5MABndWuAi89e9nhywKyWmvGhvjS0b0IkWEEP7WRautWRV7oHjvukV99zpGrnFyWPj6Mb/hBOKY
0GYZzboINfMX9KtekHw/PdMT5Rx/cLlATMGd96VJvOg2QhYWftFjcPuVPMh0Ai0JaWmhyxzNc8d4
/iIO65BQadjpWp8MPr2bDvaVjX3+Le4+wDMFSCJsI6UZupNxkDTqWXCD4CqyHUb1Hlmozk2emp89
hlsr4S6v7nQHjjXP6kLiISRa/97iHdGIlQjMPUrR147VDz9OEHBcahH/8FvnekkmtYc53Gg/tJp1
vvui9Hrg9kpAbES3jG7yJTd2hcFf4XJqBCXaa/+1ancmfzg2Y6SqA4b4H0kjF8C5zAlbNcM7CkNE
0wO77jdcA787t1i7IJFBZSthqqSI642DdTooiKz3Oci+9kMDVry5nnonSvwM+mRgPDKVxRwgwJs/
XSAzFCAFU34st132sOcC56zGB3IgEcEoz3dy7gcMFN30YasBTo5Z3GrtZhZEv3rsdM9BVGOYDBlD
VpeMcw/j5L1issPkg7RSuyv5YDWrnvGMOGwPNL1yLl7nfS/7i5JR0tpV2GdzXazwm+qHnHHJLPQx
N1TgunfviOm0eWN3SWEeQDSbMNRkYq3aFP5RAEnTdaPY8T1Fs38GUWHh0nTVOYSRDtNRnrRXQp6l
mTEIa5SKoOv6iH3odjt1rX/cONi19oW2CRKv3Zd7fYzxNFV6Xq1I4HicZuPWXoH7SqpdbNbySneK
A+Y00JEetPafN4BKoh3e96n1WZH14Fw2dnaY1YoHHVfM8a4yue7P876WVhJVsYPKgj+uwP7bxSLP
H6TgDebISyvad2IAgCadXhIqCYRLiHsNywno4K9u/G9VLtyPDaavTOR7+lYypka6rELKL6kXbrL8
XlL/9dVN8bbx2iY9dWPFuYt3KLhqdaNLafn3VfkNERg0ypWPWejIKELuj5JwN6N8q5HFZrhIJDX8
/8l3P0k1gntRnZSQU/puyBJopQ3LUTOZ0c3wQ8iU2+AzrFD5/NIP2rf9iJKeIsnvXrpiQeR1iakL
TYTpORo2S84rIekcK7m8k47Gjyyb1Siij9GkPHHcUo8W9R/YdJGeO67vGb5UjLkl+VpG4ZfJOSzp
Qv7jqQ40+jab3b9eTneMk/2cVrw5Ayu/tOxknP+tF0V4Q8kNNNouWBWXynQez8hqGww/jDAiiyc6
Z0dd9wJdOgJdKn96OoJ6KNu/O2J+e/niimjLdLepc1pj9SoXXxfygqoVb9e5LBCeoYmLBKGbg9VL
4R19cD9ETyYo6/mrMAhTtBVGIMULZ7lXJGJw4+tDtfAcMbsrFlSsvDGOhsNxO4r24K/dVlEvXwBW
VMA3AbiT39ObP1lRHLW6rxad0QCbcI4bc0oAjTovb4OLlAb/t5FWopurSgrnhFw/l4mOKmBmL5SE
FSNh0DCM/3gSNlBbd9d3Qj/OEXxrVevJwdyH8kK6BxgaMjmHrUW8jDYbmMCeZEXfOJM5enc8JXaW
AhnQ+UHkOPx0tAd5+7RdQUNsu0sjj1E4TEGG77Q38DB5pBUM/cxktrzF0bdDJSHMqz5y1qqnJAl0
Qk9gvlC/0/ikuBssfoCH1OppAifuB/tkzxUZFyLiWEOeL8dW97Lz01rmfEx9EgzRbKcKy/t5SlcG
AR1L/s51fwRfcQm6Yd7TXnaYFeXvGPQQmhqTsFl/pqMWc+KdhzsAYA3QDNLK58tv/1ydnAigDzjp
mTCUMYT1xrZedh3zh5aewwQ2/3HKSi8PLwTWNm+RIKqOyiJ0R7g/hcKSY71yDOx+6sUVzSWpjuKK
YTlUhZ/HKIxRaErZE3hbN84VvgQ8ixLObMHkZIBa7oACvg1wtwSP1CdY7WfKptzfOFgOrZr9uxlM
VNpnuUfnD8D0Ythb1qBWFuYHWqTKngPdEPVNjgtQvJhlC9MwsagG7RYzg49hSL3mDeSsbJI5RvCF
8oL09gXm6X5lOzeJnMsST392/ftQqBN8lB/cMnUGe/GfjJtuSCnRH9H2ntVqGeXPkSv17k9bZZLY
1Lv0XgHxXnSZvzGzKF1g5gzEmC7cl4lTZaf+4EnEbOpEU3Sap2NuxjsUjB9skmU3SsUaoSxfGAtm
4mcpW+5xHJXGlnarXLbKyjitMwW403k2HrEn8so+7NcZEFDh1Y9hgA9Ltfl96cnj5zcU0kLGHv07
/Cf20Vf6I6gwcPzHhkjXXXhkZHc0wxyJfTaHvrlMhrVgapgY9XcxbHBQ8ma3BtJy97ioP2Paap/4
+igs2QBQa4DZXYetg5wBCREEKr3l7sR3xFRUCpR0sGCIUELweQUM8ggb5v9gcRoUZnRDavGflSiC
milGDOutLwljNpH7yTi0AoTECaY7uV4GUs9WFxCLkqnBVNDoonksJnATPg/ZSoEfd8LfmrIS72SP
4h2Z4EbQ9te71Aa6aKtnZsw0K3d8vRj6zIplqqN53Mxq20JlAG5SJOQh4BwzDPAsla1U34l11FYF
PjtgHi04ZrgMzeKbTuVHrKOQABM7mNpxwoNmCipRBsiNce2zLetqtym5RLR+Rjt2zfxlERz5WIZ1
2YhopmDdYNcC4apa92TwoY/DaHFbJBjM1kz77QI9dyTeaRDjqrQqrBu/sARnSTwbt276EJ9Eiog9
Q0Dsr/SjiTJ6ZtBq4vBcwy+ge2UCOo6wY95wp6RubRmQ/aOZFzV0krweeAslfEd8dYN5F0+nqOGJ
BwKEP5huSbg80OVvfN5Rr+IQD+3tVpJ7OKPbfZA/XkQtZZeyYFNnbP54nMCUQdXYud4iR5XVbyfj
S37nQRK2FBbhAjtGE9vlYoEdutDIoUhKjY9+j3JRNY7m86kT0FF3EYUsvOvnf9i3LeEf4MLBvqsa
AQnzOMDddtOdKYDDKb5aX/njzeE5urBBbc0RB3gc+rzRlxiAK0rmrMfHJMClPoOZSD2e/Pt52euP
YnrjHGlVrrb6A2jiuZmaG/nCi1i6pVLSwMGl/fu0NjKT8Cv+CO3yvCdJZFqeQo3tIoWB0+3PmxGT
aLWKuaAWsrqYxDKeuU7X/D+0vGKFoWuWijryJMDyTm61+KbLegyizDa+hnKQUt5BQQT3oalynpTD
VAUP10fh9lcyt6Xb1zJ+LoCy7yE+deZRiaFcU29dQMKocoBnol74zOiNFymc5EwlPKo035/SPtsH
MChtB6AE/puTa0Tzp4Bp6AvsX6jT5Lu/kmWKCAdLiKNgYIhPo+jyHIs1icYrjGsHib5SC4kJilg2
a70xIvFkGKj+CphgJffwsJjSHlqP2h0Z+nEL9TL3Y7pwZSVmA/xAIAiLMJOqBHpGJL7/mwoXdhFv
EfuY1uz8sofnTItITIiCsrUzisQE/Mw0zZ0nzZqpw7pkQABs/tOKEoSZ7OGaMs6fpXQHabuROo/z
i7UFLG7MyCwddtVNbWI3oftApQpHR+PKqIaM/0ZWs0aojgzJLZq9LkGNx0k1oRGriuI+vZmX3YTw
VLMhoshsNwLPGNZNo7M0wimgoJwMETQ48ZqGVDfZHDmzlHoINISGxWCAxypqJ1sK9NN6S0fz8tCJ
8fkN36T1HhJBFU6p7zqMjsmgNeKVtG8peTxI/q9pCW3Dx5Rpf9L9K/ErIAauRMeXpIFYU8sjsRFQ
1SU1RLV7cHnzWtBrUwy/PbgnXNGwKGKvmd8Z/Dh8D1zZ7HNTo8Ngd7nurXIXjEb75ZSJixgS0tg1
9SOk1hgrVkQeTdS/eS97pS8Id8wBHOaIyHPEOuJfNHb/igwclTU3DwbPSkhF4S+pzVXzT7F+R7pq
klHTj07nobLuJftIitf2w7byFrl0PbG/VvYfyyjbxSCCPDlLmNr95yElJTJ0iICd022EoF0Pzeqb
S6ZEjBorVN1XGPYTU/qXjcJu8SsDbHlDUkbVcYE707qy5qTFO45Q1Wvfzp/qC1vYbL0FQr3Kxlp/
paELm/iDJN8Dgt9SZ9z9b1CDiyprmHRb3bse5f4Vl2+3jjiV3NIKU/krbGlP+TtimSs2H3B3vC43
Ofp+vVkwiSGFu2uvYSTB53aMItoXQ7xY9obHqUQbOnwf2zOV2VJwea0PFtBJQpWHOIgTripPc37r
VzseIy3JQbe5l6UppqXyazCi0cT2YppVtkuunr+Jur/lqXmTArGhvTl9pgUXEkDq1v/QIlqb4O2h
3vN9Nfwl6XDiN6cKf38FX2yML2HjUClnswTypo3GPISI3yJ4sF72sZgV4f/qLN7Pj9nA/4VjREh9
MFsrGEzcTbQ5sRzRQi0YiuiEkMHwV/qWCBPZFKoKt/yEZdjGFTS4Lar6vBqYFOqoWm15H3xk9Fur
CF7jJ6r28BB3TpewlgRsBGnoLCZJxRj5uqgR+VVB5cnvLfXRNrRKyTTFOESkW1Jx8gpEqOWBcqsf
SMFTLYuqqrb/gFEEUttMIIM4yU0MQ7z2iwlzzdXlhDqGSjPa8lrf7P22bG865qfEqMeQehd5k69H
p5vMtdwf3vGQA7xNpkmkmyFc1eHTiDJwLXA15VxCaXXfKNfB0lRCFfglU7wXiL/htHjsWuV2ZBxe
6zaz1HgxK4Nfxk6viI4YK2hbYHlkz07fTcUTc0ErwRP++rT/4bfZ14ITExnUo3pw3Pn7NbTXvPc4
1UKTAzXrP7FLt/DxgkI/3GLAL+PvUYcCTMKMCP6PIdCqZH7Vssc6WTjpGu4LzU85kSOJBe+LJPmB
wD+UdstrG69lDhqcRCiK/HgtNVkwcmaDlVoA77kyj2E8bNFmSfXDDO8ABO/NVSbdmifsRyXg9FCh
EKEEDljQYuxerHT5bb2cBxZROnIt4QPtiu5Wc277RBHDnMlSot8ay80g0pQE0HRE8vzY4g+lSjOM
C4qF5SaDLyYnVyb/hB2lnwLICWoVMOtOUFx+PW91rItgfDgo2P6t4EH5WIsOIWLLkoejh+ItGzyv
FOvbfvVyEdKC6N7E5SIbE1vWj7CGnlaY1elV3fbKHRr9griiXhM/qMiYZtH7SJs7eTBV0sNcjV0A
Akwmh4dvShU0XDws8gqTeQRpZWLbybxa+iLa6MKHLOgkqnUKREGGZX9EOsNWTj3GFsN/0kRXsJkE
3kxw5ME65MDf8pjL/aRgJXHHuDVeMrxSdKl2qJakRvLxeGJIM4dv86m8JxU0a/HWMNIVypZuX1Oe
P8AucFmYI7xowKRy0mYOdmVcs2kcJnX17+ZGfWD+3xM9xLAwAxj8Wj8cuGKbsVGyGRfOKaLj5bz3
0gEehCzQBY/MMRv1AaXzhKEnpc5dm3gGZeJyCz8faZ6Dcgn0erXzqsnI/A9WVZymADhAW0ERFJJ+
sw0q5sMr9jqrRiLDcFSK3jZoJKAnO7pegKNAJFMp+P1X6vGAvc0De8fUjkrJUJe14ABcTTQTzhpY
T3xALPcsprXLoyqTrRb6GbSF6UbWHXyBpYnirHspkXgwFd2YEDzuE5GvihMfWdHQP1nZn7TlpHF1
mUi9Q7obg4s8kqvFVXD6CZPkeactXV7nwas+qI5pKWfQ8ggEBeVxkQlSm+I9o/AfBXDvZYqjpN9g
WYnqC2iuXmOTpAh4CeAeVqdmn/9H/aCbRwd5GHSizM5pWutMHr9tHZvTMFnRjKzO8MVCRe6OykRW
iwB4XrtMjNqLna9TIzJEiAzpNpgVXGNpunaJqVY0J45IN08dhfVNBeKWv/yn3lWBNAUQlV2vMLD7
gc7sMaH6JbfQwH5RfjmXkKXdX1Qb2suVR5+jYqQyck8Z53i+Cc9X5z6pgTLDvY3gi0BwewtUYuxh
WYfATMZhO0qIcZkAEHwSYhIGzPLVknx2U8a5htiwbRkNr1ciKG3b1pbvEa7jhmlZY6tL77vjsvD4
C4Gq9l2RP5fWohhH4OBBvFtUvkwBj8iF8rXtFedWwQlox5/qeOdz+9uT5twAEu7b+/fpzsHdac3w
ZOS5J2ELUEUyrvq8prRGqTHXRYVi3FCJY2OKkMNvTi5gfo/k8jhNBHsq6oWIZ4jlX9ztVBiclOuq
ox1IMqDCzHyJLbzMeV9Cr9TMls2E1qkJLfteE1WT/hU+UpfEJfaECoPT44jBYOz4S5p85MSXVwWT
kTKlWPpqVmRWAFxdnMg4UbqqUWRO3rkMBREdm7KuQ1ldrtGlQl09jeZePASUv6hdovJge3XGVehr
2fxaV2g/aF0mS0Miwy3A/7Yem8Vc6V1CM+bVr/86gflUU7hP0knTU4RyLa5ipELvJ/WHNDSc0c9I
uI9O+u/wTnAF6tW5suTSjkdHqZTBmtgw55N3haIgIbqsYCVjXrcwRbT316gN3r6m6gX0MZTiQqWV
A1Lh3z0ws5a+s1cd5x77hA0BYZyCn4qtIFczcG8IkS8bTZq3Wwupnu4vDVutu6+rqL9XI5AZISHk
S7GlotncxPsNJh7OeT/nfHw4Mz28xR2INU1qK5L/m9wKSkfH0jA9JerogeOPzHJ7Nh8IZNPNlkt9
131QVI1uQ4TW2Zf0ev4mKoLB6GEcPdQ7NjXvii4bIDSNUevC1QYov7HYkcEAGxPu0TpgLgxQxCj+
jkavNO4UoEmVx/68BwCN4PiWEFBsWHgKHfUY8TG6KTiZuKdpG5vvU9ptzGsL87libgZeVVNuMs8A
SCDrcQ9KvZg47MXLGhxYyx3aSV2xW2eKWA2lgQ8r58A4S9p5SJBdIt+z2+hALqWS6i894H6hfQ1e
nir+T0lzNk9xqB5VlYYtzIjpScVaGVHcHq9/IG1SJ+qWocQPcWj83OzPID0TJt169bnzOtHB8quX
W+RnrFo6Q25trAWEI5R+zqY7X/QZVpFeAzP0VpkQxSwMsDt4qdB2aNNA7+ONOA/SJRCVn67kNpkY
xLRIf98BGf2eEWfWWOMYMZgzHOQSEdtBmQPiJ+eJlEfNsXpXPs0D4iJOub5JNqI3VjEJmWSKc1T3
VfD7V1IjKd4SNJEvy8FDNAIPPL3DLEaCKaLtM+HjSP/5rYAA0+4ynWNug68iodN/2QIFdj/adZSQ
fJRQ1X2c25ULSBsEtk7oaROvw/4QUu170jGQJI433Wzi39p2LOSHCyG7PjC2+3WUUk7oDaSf5nYf
peqaPdTCzYa3Wly0kkkaWF/WBYQvL1wocEDKHLqhg9uPQ0F9LsxcimCrFGTzSRXmeXZ5n3MCCvqE
G4NiFmZ4XsqYG5fnAfTOXKLabxY3kRrWoWkg8wj91ZGaH8pnytuu3YzaO4S3h22jJCjnj3pQEIXo
K3eaDzNVDC0NOYAqZsZZ0UA/Aj/IjThdZuE5Vqll1K0RRI2fu0cYC4bL4vk5Gnh9QcGbBfdaeOIX
VIQALlslO3dVWEpU3J6SOHjYCtrKQGf/CQMThXC95ilalkIkO/ugxntYOeKYBucCre1oofaLZKDx
ZnwJsR3Kq3ppvTdLQ3CmuZYz8Opt3/YGtRubwb1HWMoJ3n8LtStj56l2trBmozaffIE76oesdsZp
oPYyOzrhQpeG9G0iQ3UV0Seu+bvMOs6tCo0OSl80tJFODtJVJ+yEaKa63LCV0aflnu9xs0eTqjhJ
1ngcvDkFP3uhNuQjvToHUMQZtMDcccaD9tuu4XRqbNd57iAUoXiwDPhuROl8UgzkgTHcnItDzZMW
Z2ZwdgWYJS0CrxxOf+BiIJYU0lEF8/Uh2xl3HieBDQxMSTvSHzUn5EZtD5c/wJDBVj8KAy3arr4v
q9T0vKyJ7S8y3KUKAX7dD9GxXzSTAWC0MevdbNzsoM1C8aKPDx8ar8S635t+tdcjgSWo1wi+WLrh
WXeVH4C3TGSbYEWSG/GDCIh/RDaahfXar10GMeZ9FqSy97IfehRlHjjS22+4vnZ0vmHCwaxEa9F3
t7kPOXedkOIYbs/mWT5mZhoP/gkQR0vZo5JWIe52vRVUfk9yiu45IlOvYTn0rmz29Gk++AXuKHQN
fOT5wsCSH4U1ITUBPSzLQ5AoO4zQJii4g85ZwfD4dqj/X9eJnXSJcU6ceg+7B+vsEb9OnPNMW9Lh
dTJcyppz2XmRuvk+K2MY6hm3VHt5GM6jD3rQVbVVtySmlAJU7/GNkJVHyiHnDFX3cJZTyty+aWaQ
8eMTGCXaozACgqU11tXAXMZ2cwGwJcUFLSrsayIQz1sATA++cAqUEUUw0atSp9MEw5CPeGlgBuQl
AdSJdqXtk6D6g6CnWFWerSnVnSPpY8aGAMaJHFd28IKeeSrNtn37HT99FOE/T9h8Eg4sqaMoTkz2
ag2mqLQA1s0d7zdsWbrfDvKwtR8mRxlZuJWuW8QEM0BrJd8Ii6lWKxf1Rjz/zez4e8C00Q7mQ3v+
yOU6Iuw6DsPGC8lR1uyRApSiwU2lixhIeATW9ChoVs2ts9rKdNggUCLmLIIqcEdT0Wre90VpKUkA
FSRNMlnqNiBteuO1VTGTSRUejZTjRl3aUzVZ5/5XN3rOEadEXe1wbBi4ddBXqwmgDoMA6iBgE0YS
kwgFh+Iz4v1ue4dYlJzyfYaoAQPYE0/ekdarS7tP1JB6amiMcZfpf87F1eXDiBblmgZlCv77irqz
veFW0F5bmvmTM0QI3OC1errMX86OH2iG0uM1Y+PUr7jDakKdA5Pvpy58Q4U6THGiy2+vN2DXZEuz
1uTiygvg0h5YTD+Dfb2H3TxzqctM4byS8IFUqcVzGaMuSXlsJMb1fu/1zdoFA6OZRmQqoseIVwI8
rMEEin03hHFbcH8vkEckGHTu5sLHB/2rmyNbDcwha+6qctU8ZBuy9i4EsSo7Fg821ghBID62Gm+H
Z0ZLVQMb++HEQLXVPeHeXM5eTem5XIbmkS9njBxQG0hhxdNXxuFSMBYehJQc9W0f8+THES2Ou01Y
tn7+KV7vFnz/UXRIR37mhLFSnIntnxZHtaK4r1M//GE1cHiCnbYCktqjabeVxjV+LLX2/7VpqWKJ
CbfQlabBjb6ClSG1dATiyj9SXgTD9Cxi8evZFzJvvoAPQ6cuDUxyYBQ2/Bqwr4nCxFFtOtvPDxx+
okD+YefpTAk+g2JWXuwmZtJuCcqpb3DlcHnHWAtD5F5KNng9PMd8Zgwem3cR1C6I+6L2Lf3STQvf
y2DLz7OUGFY08lMZ9K3bon5LyZJM7kjDDHek7w5qifCPMGJ+JkNMn1xzK5IaQ+BuoCcYPc5Kuvky
Ag3hoFJWYguHAFoG5ZX9V3EkyBXroe1oK2LYM048H9Coe2dsNub+wQIqvyC/oDUm/jIhqcSWz4u8
HyYStQF5Qi4swndnwMnboRbb4GoCJLknuqjmF5p0Cg7xJRXvsJPyiIdAL3VC6/GTuT4MjpDJo000
+28zawLeUpT3W4HMxF+4KisQXfA+bdzC6J+AIZ98Xext4ndZymSNF7Qw3Sg7gQ6q7Fbrk6KgurbW
/gfjMSFJvonqUe6aoEc0sMmv2nHNuyH8BoqGWis3d0oFXdahHWlH5IbBAn11CimpfuJforVPmLD+
hshLI6SIY6dCszcpjGAm1+scZQvfj6ubfEw2Hm/iAqp70OLSVGEGvfkwW1WFPxNoGE/XvXU572si
csVv4L5Vv/WCMYy8kHPZXL0oophuNSISjUjTTeyGweEWZCGQalvf9zoVR6NYfOr0OX0vVjcV9SYX
zkisLnE/2MCIb/DZkIuEeKXo82cVscty3Sfi9Uk2m1J9w2auuSNDpkA0zS2n2cPBi1Gt3OLEiHTu
+rNc6orehBcPfH4B2UXVtVdSmGzW/uNPoORiyn2UyAacGOPkJ38RnqIZPR01rR0opGLLPzJ285iG
F4pR/LoxXQ8KmVaph9+y+oRhnq/W9nil727DLd/nzUaohRqBB+slPVjvnaeVxyKVWwCNE6yvhw1S
vhY6gFdVYDgmKwqf2OfPUAPZdVkzKIBzf46Ke5HXxzjhCekaR8OL0mAJnkmFvhCfwKPA1AB5M8OK
kD9rWFnIyqd4H43wNhhmVpWfOBmOUMnypd7uLcOK0mZz2F4juTxRm6SfBpJMnyeB3mzwQXNjHxk+
i2Kk39WmQdlUsBniDF6m+V6yD8aQ8hpC6JPXDsn8H7BoWvou2CIC8Cvsb2UAYlIbHsBtwRNkKeQG
q/2ujJKXQDko2aFOQZnw686JrCdZyE92aIlGW3GfrAm2kySQktCIz52Gce0VrQzez809pSv+jrUD
tDNQmI7XINqXE6bOiv2yHR7IRhdxkb8J/EKa3rEfn9SNyxubeMDlk9XFdvryP/XSwbNqiVsCRpCf
UnBCtfkXHHtm0gFBFFovgIbQMfCy3m8d/AT2G9LAYJXzl6soCEN2wqd3aJdPDSYsrb2IkbYXNJoJ
pgQcEOGQ/r26fdAbgxGGU0uYctY9Ay5I+xf3ibe7t0KjpMmLYiMaXv1q0BtOExsQ9BG9adoC6YvW
OlLQgq8FTSZz9yg5GEDHCOOTtF2H/aGCwcR3KJ+EQ0yJdNhZGBqXHR9QctQGKD1ufncIc0mPcIg8
YoKSid3dgYVKngkmQ/inJKZA7Bs+e10A2Vju6G0CvXRTS/+SNJYImzVa2dBfI2kA5o4XC6eh+Ip4
EVISu5oCSb2aczCqZICUiuXx+d8it2b9HPX+uzLVypiG6wwMZwy0/Xh3mYWJtmq4OUzccvmJ1GxG
EMhoO/IbAJEHWwrEjtQvzCG2itYCd7Z5bHXOkfJtWMu2vCmKP+yXNiJ2uoinwYH9hoNyw27Ks9CL
uncyeXqWmhr/IDootoFAnpwmNoSleWVpAz7u9c8SwGHfd8M+j8AxbrEWLiPc2XmntQYMz/uyIVmR
/OqthcHr2ZoEjtaxfa/PnHsZx11MkOWgoKUgP7pUwu8AxAA4igTqvQz3/D3TK+OZlPIKxiRv1izu
hI2HIc7cW+jiB/g1fYXs/XQ9Id8sazwPujtAVEp80OhSE8nhNqNkU2kn3q5hMSZMfm9gG6Z59ZPz
xMmQpZXoPS3LCdMa8tKwwnFaLH3mUf8e5NsGD7zGYLgiM0jFra2wl+vlSIK5gTjkMvSxRkQ6j0/3
Otg8ybusoHlX36l2NECNcsyi1Y8Km6Z3/afs1p0gHv5GpT+0guG7ovIOE7UXxZi+0aEe4JyI48BU
foRtroJRBwzb0KNotX/LtcT/OkzjcxiAD/MyN/95gBjjifVvs+4uijgp1vC+f7+jWrGheNlpqDgh
UsVTENjbSdayoRML9MNx9vIJTlVeqwXhnLrDoOuzNPWhgC0mk79qXevvf46c9JfIiQz1BGKZtowd
fKavot9UiMisk2KbwPhzkLNAQU5B5Nms15y87l00vXB8Xiuih68Wj1gqI4cxMkPNk/kaAc3w/Mkp
tnatbA7721hXu9LHMmU8TRtajBb5LVcFcrPUmuoHuaENC6U7KlDuGtrsneI8pzwgZL089tYeMBmV
dBC1Ba1xSfoq7BVh9DOGD6zmKtXPBZ8LruIaA7d0DLzcBjKulPssM1irtoQ66upCIyVboKgagEc2
3MWdr/bV64ULRDFXUKwj64ZA+fLNwarGw9aVsNXUEZYWn4/j2Vfvfycb7N4Xar0riYP8snHzuG5h
bmX1FdoeKWZ3AT9VTqf3Zs36HVBUThqeKP3AEOtKwCsxd0aHJ/vUfiYK56qW8k+EQegGTD573PRs
E4bvP2Dfy9caGDEsF9ZOEv3NM6yCATD3Bp9GqjgxnOQgZMWPLCison0ZAJBsbKjGuu+OppXUlFMG
d8aUodNxkP8hRap4R5GjFLt7Ejvh3IyDmD/gnyB0e+5bn3/hcrmKFTZ5PxkBCWP5l5kCpgZ82azl
CrzPRHXg6UEF+Rb6Y4yXlQfpMcpjibRsM/pq+Ke5CsBkN8/NMzW1J+eJ2uH+d3/tg9Pam/aFAU0y
Ued5+o8kUMjK//pF7WKubV0bhAs61VbXm7jnj9WnnIwlkyfsXklYczxVK4gFzPMOpusOyHAUwSM3
lbvV9THprXswj2EH0G2xrdzGPY0KBA9hY0+zwuyeRQWPI+qGjIcqVvWiNYHZAkf0imWi/N8gX1IK
g/ymDpNXcXrWUbo+c+S2ovSLX84fy3WBilzkjQyupgTRNifcU07gidrdTuj8I7Idf9unecX8saHR
wCo9ukMKsdKgapzY1dbTsOl9onXWaGUFg7fe/58AqHmtf3+zAM03HILvHWZ065vAEVjG/1Mrqpod
5SMiuhegD+rlpUUJ20mhubLSREOyXhbjDKBN73sElPTrGZlBxrOAfLhZW8E8hkSDkP8Em7qdHnjl
ZuKuLrjP7/yZFpE5zk/4deotTHC0+v0H60gHQtrA+QmwFuiraTcT2G0WOrR1FUMEJKsCq8aCZjRU
DlS8IvcEdRcGDbaTdtamBZGLBJl+GpCr8NsW633I4dZz4qlcL1irdQrR/nztDjUT6DZqHIMXh9/A
T7RnxQNf3F5auFdvkzlJRg/nqSNUPst/PYs4DnKpQUley6uMNFFe9bG2sALB7XqyfCJod6dRIlnU
VZMt53VbjlZL6tCYPEouHi0mbYCV/dE/zrSZugxzHqozH6w/jbzOn8Dnaq0koerzJ7CJXO4eMNPc
nck61bf9vZgijLZ0CsuonUcb++zvruYESCF0lYpzj8f261ADchbEXGimap+ShkeD116lHXawU4TS
doDRuHh9kkEbAbWoI0Kpr5/EX5eOStSSjQ1J5zGmvthu9Bol1ipVc6xlGN2mQBk29h/dfnEEmFf4
0+4wbfqnT/epoO1aq80VqfBxzMa7TwzBCBBgr0bKB97i3zHLpKSJq3pookuwSLIYVkiEsjDDhctB
VgzqsS8LLhUl5cTSRDsY1ObH9j4YuYXn5LvW4m6IbHVTUSeFze9c2Fdve6iXqmkIaIsXX89YE8++
3liqmqi09sT8PEu0+tNRUvNTT3XxjWnbZ4MmzR041CtmlQp8Z3VdLuvvFpiH+qqyADH2/Rov2+vc
vtasQ10FZHYDOKgfTxyq565qW73anYcppJ9DEdin6k1lzXj58R+IpHJQU7iHzEXPSZpae8Guwpks
3L1XJlH6OhCnaDIC1iEx1aJVE10CMbACtDBAq7ctHgpRhBWFpo/yf2zlMpuhxA4VVY3wFXQ5SH3R
4YY6+6ftjkGFyJ45j7kDz7yKTjHXfniMJIkMniBXK1CFdS5vXPtwDh3MV/4b5GwT1SwtemH5oKX3
DTtYqHXYNXADc1ug84KGObMxPIF+9ISDdAOnNOfK/sSc69zeWowKT7/phqRlX+2vFKhiL3W7QnpY
XoPD1V8v9FJmBLgOgAX/2ynBc3ZExsrfKSwPmiUxuFilKcddtIO5BMm+DZME/A0JZAoUbzMfwrOA
Hj1Gc63aV+kkNaE6peu/b9AKhL0C1VLViXQdQi2dbkfQdPotTZbulYdAzxQ9zXS9I0JEz6UCuXe8
sgQB+WKS/2BHmlP/srkEmYVhon3uiBJ0iVCQZ9/Spieq3gCed4eRrrqZkcbSbSfapanHQ0+bEjIG
wiQVS9uXoQmi31e/9YbyOJcmYOZs03KPqDrUq+8+KG/lhyQBgolRXQUGoxHgkai4JtB6vabtecme
olgBEkXhCaKdpd8qJ8UIxptiAdleRTthXlI7jzvTvubl0b9SGbg3ohwbDCmSea5UvWKEOGTUN3qT
V2CJAK4x3qkP77npH7yfO2PhZPQZr1zZElWcJqmtFiI50JASmem/eb/Oy3svZ+46zUn0b4vVsMPj
yuS+DK8p3QTgiz4LT5vn+1CnQMK01SgSDSdZVP6lts45Qeb3mfGFwDX6HZ6UBI290ZyDUiNbbkZP
73+9laM+XlEl0fzkNfqhUFLeJYN2USc5tZEzpccZJYEVftP2ZdfTTjIePbbzMS1T4ZM1lGsnuaTK
l/hhYyXvs/CXFUnzK9FDJV+Bnr8pAcgmWjMn1iq7RX2WMfwl2Hn8pqQoGW5rmnMPClsmsGilPpdg
XHbBZ/tFgITBdKCQlnRZEPD7gLCXFPJchpFa5yBrJpk1Al1GA35dinzYD2gaMPosWYYyNdL1TlSd
eoroLnWYjT+iIxqk5HX7KR+L5PhlJYnlBQmjtCjzI80Kf1cLTz7hxDbKZI4/+rrAcU84ozrVXbwE
OYaNpBhOUB41Qzbpkn0Y1bPiWBis/SxlLADuONd4zoNLsdG+/ImKvxabjwtYGv24fMl6VdSs08nG
ChErvXAbe3KX9AN5yzLjJz8B9bC5HTKlg++8gIc1urY8FkCTdbPdfAK/6sNVgZfPtuDf7SjqLGMw
HHtr2tkt7+gA36tDZ6R7WNH6dG1gUdLXhsIyoaEPZhzyVwOtGfxUQzuod7J8YBhEwlbngrjgtasy
nFno8wBp8GFQ69EW/2T0ETnTNVqS6VNuYv/8YX5OQE+AvXYU3uOEoAJRvnuRHPxp21DS/0os/MfX
LTUr6oOcXIioYPztXxBH0e0PmsCdWvq92yXGNQXWOK/wK6emDJSPwi+Ekzg930ma9zy4QBEKmbBa
ee0WjGXSOoZq2DUjJhj7PtVkoBAnRTLFzjkI+YsrqprqKZAgnL4aSdC1DJKam3EV8R4SxycV5u4n
JtNvT0n+RQvMGbTthG+uRe/fz1RHy2beSmTUC/BNnwYy3B1mYnfcXhsh4ISN71Sa3nnZYqWnHAHy
w0OComs625iKUpKMKVPewbHhlA36ygHY8n7I15G84gTzQgGz9tVH0f+zQmU0/qlaJ/wolK931YX2
jAJv2bZ1XbtipM8Y9VHb+5pohGZwJBwxnmTQx/cPp9Cj356CglLR3Ridx3c/0MTnhAug/ymAH/3O
hGKCm8ODC3JVLj2qDmYYKfjfmfgIPwVH9kMC4/sY7EMskGkwBWgzEgVJ/qGtJ/uethp3Blc+lE31
wvbxyu8BKYRxrCmXW5sUXaxINa8JgRgwkhUdIv+6lOMYh1I28Q3+XjG7o7AcVvfdYpVk5MDunPPv
N6U9CjEh5Eu4Fz5pNIGSUJiTHJ/07M5nXtwbv8K/icGdtwhxCpygmkq5Y7tX7P9jMd9aT/Ev8v77
g6a8c2V2J6t1Q+iSnKR3gcVDGLyZazNRvXSMd3EpU6HVSSFESYV0gg06fzeDVkfVoaNwacr8hvnn
WtWhCuhwIh0+CvPQ4flg0WAETD3HHgtdIqc7KmCAarm29y5maLk+MoTaP+bDIK7Rs64BCcdB3aVG
3t9sHp+Xbg3gRvEa/38ke/3TU9f4OfvEDNt9NKUbt3UizJ2Ix5ippKc7DJmgJCCPnCZZt/qQVbrS
80alR/zd02rDEUWGYS9wJsz5nUMIGZ7mvlzG+WgmAF3D/OCjvq1dIIc9id1rncKz370+SOuZSyxy
F+BZqo7IlbS3ppXw4hVtvYeutFEDsxMka9Luneye38iuzGv+NnnSxxjknXagrzGmz0eAgHzymOrZ
RjV/oi+JXMdCD7wnxz+bTz4S+MvZEQgF96zMJXcFWAzpuw7UcVY1WgAlLMyhGanWJW8ZXoizyNTY
jmyY248v1DEfVf8CiMkchGCcrR9Ll8tmsW9jHHRzn1oijsVpK+4TV00c/0jfrAvgiOArs9+CH8BC
wz0kVYE2Ue45p7oLmaEBwmJURB8DboGnU7mjodHICyKPUk6ywnTuVesQkLFd5+hK013LlFjA9QoI
A6w2/CRfj1WERrgZPDMwGGEHZG2RAUVK+irFCPLy663qspi8EdnfwRB4j80FqJXTSmJcz4/oOdBZ
Eeo+s1WR0qmJ7DsjzSGqkskpwRRxMvM71tFn2BKwe/pFs27FS+SuHsQOZrU75CAk25VOT5P0sXx9
J5U7lTFqRi9ZvbMZOwZGZnQhH3nU+cmbO5X6XqbnBvwHD4d5fEzpPuOlHcwnXS5R0aWPZQL/BcAW
zQllt1cq2TdpDOkqa4oUDSA4fWMKx9jJypfXQj4hYX2smztUA8eZ9ZB/MYeNaytYJKcc0ZsD09oh
m+1QFMpdGfIYRK1J8DuUOsY8JtkXMaCYTeLkT5HQJXnjPknK8kNO9VhEoQBdW8HOrbxTXmUfdq2Q
T98P76ILzdpzP4Q21hhv7cGvJS7t4WT3Yox/efgECHpGZykGaqMsr5MD7V4q49ia4AcsTo+esLda
6qCHmCaOmtnJX7gP80Mbiln5j+gsgWfkYCKEfuTTObwWAL/nhn8k8DMH/rm68QV3LlmXBs4LNPZ2
ZAW/kGeK7kUKNRrNxaHs5poyZsrrjMaUfF1KuLmEgSwrheP6h4mGKH6w/xpLz4TKTEC1L5l6h9ve
sVY6XQg7Jku0BLbYwLu0xvif/s6yVtm3Dt8ScextR9i3DKXlWaFMhxh5/wUskwHpnHt7/k0tnCr/
eZH3hajP9QEA0hepqTnZFSAofqT5dCnid7ZIG2qjJ9IrhRF6MHO9T+NFWgvqX2A5xvbucEaYMArt
hPYpTAoEjZK4KOJ/hlCKAW/GrT1bWnnwLxEjef6h/5X7fFFV7dR3NFLYfTe4VMo5tSjIgslr4/N+
xWuvK6HpBZZYtAcoGwdwMPmqIwOKJWijXlWv5Y9Y/VP9afrNT1zAqWc9wIxzm689QWE8EkRiYY3R
4KgI3UlXZmaLfm8gGyOep+zz/6lI1P4TplWHyj9bMJxBJNrdyT1t0rdf7OvWU/9n6MHl4FpSSToL
2wc2ER59ZpYQcbiRLcKoH1bl/f1gGOIyXM+BCCzQHEU8QmXRq7tc1tiIcFLpPx0cwHD47yFcLkyQ
83HkyzQOOkiMevi8P9TfEDl86HIDRwv6D39121Xad1VkgMB1GdDVi8UvV+wtqwPPVQK2KP/AyQ5X
+YUbuCyLdTpkkeEd/QPbxue5gFiXIDfa3LCsq8wnujshYneTfpLqWOHBlnI7PVRNzlB9iiEokxOq
E6wvhaWxfjJ2uX2jb1oH9SFKuZaSQj64opS03go8DX8SHJa3uV2Q2JgxdRtlssnSeren3imurPbk
Z0k3gchxG9nHB69l0g9p0czED76tPdMG0HZrhtHrFX9a8s/JKvngfr9mz/vyM6GR84MXFEwyQ82T
wRQG0CLiZCbc1N9ROPkYn2lRUpZf5OTxqZ2Su1PG2O1gLdJN9ONpR4F1dzwEfuffWadDNwQiO7B3
ctHX/CkXy8WEQUrjZGTCHEbePz5bpC666wzf2OzkDpn8kgKxg8blE2A6aJHdlFafZ/I6VNEVk61r
qWbPzrli9AkmmubTCE+Y1Bf9CCfz2gA6vAeN8V6k051clUa7/lzVh8xg9TJTjm/XxtLMgq5iafAw
mq313bv6bFg/EgY0SYRM9pUzW94TkSXgWSjLxVh4bsZK8FZ96e7rprb4+hVGWa8/FhyFb15gDook
7yBGiTx/Rgmv4AXD53nuRxH//P+WCju5p2mixuDywXFX9tMn0tNy7pWZpaAW3SLC/DbrK9G371dm
7JOJeDM1Izid+YvRdudyEjCwnF+blYSW9uz+a57bxIMwGFP7dWzsS540Sg/5D5lwLYnavN60ZsdK
SDa9t8hPDw4uztoSWAYgEKzJ5ThZs1TRW4/OLZJFgSyUs/omUywrZf4i/KolJUBot7HADSy0IQKL
cG7QS6rzAgcv/wBqv+XIhdKVnW/A8WTcRneL2tIg3aFqF2tirJy8XuNIBVRv3XhHJsR4qxiiWHIA
424DS8h5ZSKHBetF2WZkJ04KkJzI6s+OW8dXIhkkTY3ETXT3csAesGKz3LiEdK1Ir4egXmJ3Otkh
HY/bBqaNJb6COsRA28Vq9/G+lVi+RlxIXyCN99D11gRJlOuGX2Oypi+gcj00ah7KnxlxhTbgZ2u2
XlH7c6LPWoUdzGw0aEvIS26PSY5hG2e4Q290Bt8iTDVxipOBjtWQrepUfXiMdfPpygYiwXG3hR7Y
QQyIwUXpcchbCW/NiFAeYnDEvK17Q5/a9SMyzsPvvTH8Zd3SWO1iXxhy7FwU87iU5rJhmYD3+ezX
SfrjLPpw4hensn+G9biKtztBHmsrHkvPV10EROWTLZi9l4MkDZ4CSYCJuQtNhzkYMfCWG3L30ecL
4MmgRkzsRQ31RJ7hgU2ApBTgCis2sklygQ7XqJMc9k6O6AHIVU8z7MFuw/Pr9bmG05n3322HLSs+
FuL3U2PruSD3dUQdetErsplSmBwkhqpfTTaK9HaAkS3+0b/kaHb0To/U+FPX//RP7Tum2ofeLU7R
RDvuPDh2bQQRw05CEQRKPtdziulFR/xmuJJpTrfvr9Z2vucUvNdFhRjGmion8ppprlapW+2nsNDf
W0Uye4ZL2UJ7iNi6fbBXg0jiiGtSRIGdAPvlrqrhvzLjKIzwjT6oVoUadykOsMf5AwQwgWbZ/NAd
C+AY4evIX3BPhwMUZXFxuMQCu6iky2AGkgmoNOfIjfZSQb/cnYbEaJS+Wqlee+b8sHSoJpqokhem
1z1YMRvt4CUSY7fzTjAAsscyxTwPz7HucXZ9QMBPg83fSePB0epOxt7OPG9ELSP4G50p4KOdOwHU
c2GEx5RNMhOu6b19WK8edsRp16tgytRcVx4q+2KA1jFj65Ybb/za5Sf8KDEnBhhRRhtIdOGxg60J
Yd8BUKVp4Hshlb/3mP7S4UVs4hYyoKLMn3AkBUFKdmrSqISbZaUV+e48nwiMvlfOUMRdAtc8sEYf
B3xCn2CUAccNtTZHbTxYLQMeG2LKngR7moLGg2DfRjxV+TPPIyZrAv7CysyCmcYFPZvuhIA6t44i
/q639il3HdbdKhDGkfWW6mQ1OGylCSwL8s04AUnMzwaYHvQEsqMGlF+nZ+MM8WKgT/jww4nc7rKz
MK7mWPex8adGMcMJsrfiTRGX5hf9dXdWZT5uza0MaSCvBiBJxa2tRUOTJ2ebZMHw20lGR0XdMaRj
NB+NIYP1rTqH2h4pvc7dBEFiLU1nzwpYLlF/PyeHj22k9bWRmt6t77w7qh+6Ef0x4OgQems7ipvW
INAY26vRGwZ1Z23npIpnGfVZl8aloNt4jN9Z9RNcpyOsdrqc47k2yJvlegRw3+bMnYwgolylohl2
wFLm2qbPLtYbm6RjTV0/2s8s8myTCBfmpn+h0tSGseotGEcvT7hpSLj5ZSxsVQobsdLX0GBAVbGj
tkyB5mmqTDZmjgJGfsOXRpKs2vfdFmtBz7BcP9dtY8AuS+Utu4rgJTm7KJjilWHYf+2zcLNryNaY
BXV5yNc6RaY0/xFLO/ZcJD5M2BFjzB6HWze8iRX8h6UYn1PZDJ+KGjpK0YVTSFb4IWU6RVGdVvWj
xamdXLIOMbx6J5G37htczdHv8iGpaDgGBYdJrOodFIgTXAt7b8dfny5omGQeo6kYuMbPYXRMvXlw
HzBw13OXOjxOMdDvQKyTEtCmM07LLDN11Gc8ZMX3UvGoWguk1258+3d6RD7hSC1ECio8jvngN27/
+n6J3L2ZYU2HBXtRKblchVNWD1sJucOk7FMiyyUvdVLgJynSrhGwFrYyl3zL4SJHajcYmAcd7aoe
SzitCidhFni1ge9z/n/Yv/VOkCCcafATwS8YDQrdt0Hv3IlewO8DqrcxgjxR8PfEmrQxzGmTwxim
zm3cQ3BktZjLIQ8IA5VldAyL0xiLhmbRF+Fy8e6MP9XnWWdCyLTlPAbZGxayijAgzgvvwFwpuzdE
IG4wd+LLjzx2wrjZ9x/5o+UiW9RTU2oIdJIGkS+OtOOFnOjQ1mIcLOmALuPG7MAQXsHzg8L6OLca
KAesGXLh1DZhCROp11Yx2n7Q5uXczW4T+o4EEbFEFV60Vlu/bkfu2y9ATiLUlVvUKI5j1wdEI2f8
EORh9UBrsoO6fJDglfQyZgjp8USFA4lU8QbCipsPx48fAO6etc+FFTDtTESjaWSv+aQYiHcOaaJH
WpVF1jUtsleu6Xt8QI3+bvtOweqlNgE2nde5Kg5FML6muoh17SdKzyETL02C4wnwxorGFkjxR2sG
YLb5ZKrNQjpVjuY2rtWisO7uy3K48QTYVCqlMeoWPtpzLpf+wys1Nf59uBJBPaHTc6R55UqCbPz5
htSZLjmKeZQKj2hjOPncCfh+bfoh/wFGPCpumUI92trz4S2qfCYHS8XLgfC61xWwPswfWGBy1yVb
rmFM236oE3cT4daxiPyI1vV//yWmTOrIbl8jOgXZO4+gj2sLPprEKDsr41cb4NgRIxLBWV/cK0OZ
YJM9Lzzt4xFCE6p2r6WG2W9mW4X9c6tAfnxOi3Tc7mZAXGdT6CUmwRvJlvpsch9sNCXXuiiWe07A
HadUc3GiV2Aq12ocQFlm0xJH7Pm6HqGOYXxFAOs99sAld6I0578zEuiFne3Os4ZTHOWZaOjcnHJ1
fYVOPBywZFzajHPlNl9uJRKQGMWD1EiMWQXZvTjrQunBccYjK7dzB8m7OPJ5byqPBBqAFS26rhRT
8ubVoY1uv736qILjKqDxdsjCMZXxUikeZm9ICsDa111GD/ue0n7aXlfJCsm5s5hydsfssfGpeQMY
Zf0f+5qF+cVPGE/R6Eh+FNBmnPlAXnGmdtCLMtvUbr1sJqMUCbbPvpk6ImojlMVHwObtVqLjBGYQ
A9X5cjl8OAKvGKtibTzW0wRGaOEyMHymPe+L6cDybgig2M440s1ZBn9Kggp7LcSp2AEgFGleuEuh
z0cnG1RHQBUIb+dxxkjF3FDV8LSyF7bg8ZyK+mRMSR5Av/fh7zJmSrGx8uu069siv4zwE3C6FYAD
mDyjyggBnKwFTa/cy6xTHEy4PkxWgyuwvwT+ruycAJ/0fQTC5ZLwsi4mxF4APT5oB4MVvctbwhNx
al5md689E6kFOkDhYwlyCFZMm8YCdWBeU86wV57NV6usocw8Z7B2tVgYYu0+I8mlIiSRA/ax3Cro
l//mZ42JgOIr2QMjfM1r7x/hfQcN7GZGU1Vn0Jd3N/UuOfN95w28ygwNor3cw8zGCNbW6D/1n50w
IFmunfsa1jBpplJv7PQM3uTlS/GVqX71PBEw6P4vJm+2GL1hPCqaMez4/l27foavyInYCcORs7/p
0rxP5MZ8ln24z/epVyjy9aeWZ8pex2u2k0WVRxpUHslUG1EAWmdCTJCneXXQSQR0WHnZXhoRCHr6
5AhWIPBpRAFFRyXXBd5W7VfLErhOAzHMe98vef58M/8iLI0Jf6M+Vm5BwXvbfZvRNVkUqu/24oQp
5/VMvF61FFCO6Yf2fESc91JcS+ZoG9+6RImaHSdSvMneddXb5DSXHLEoinnpZ/CXmSfxZ2krp972
I7f2EW8292Qwlyc9BbbGiSpUECQja8cwRSxWFFACxOAxJEEpGB+m8L0z0gtnfopgvrPweW0fCKJp
4QQKU+ul3E94K1r9oeJV21w2b8+NecWTVWSNqdptE1Aq07wmHcuCd+HW2vzZRgGTglNCAXC4yzog
8ql/0t9+qdW+xUwl77durQtM4Y/w6N01LF6KOMVqtoYqtv7YIpdMuvopuB9kXmT3VWg9il0mRzq8
XLG1ScfbulLhf+ZUu3fn2XKOStqdzANi8wBX2gVYyUKrdxJS9Y/ciMo/AQpTd/hUkaNzxW5ZU91Q
QnxGfwJTNxtci61C4nHhr1J/880nhiN7lueOp+V7Yo+IPOfAWqZ6r0+BHMN1aYUtcwQdvk8UX7Xm
DqAWRoICc9WqTD3M7z/cOgQB7mt6Eidy0nItMsElNul3IP1T82LJxP/SWmdAe5GfKh0iAg0NTL/g
Aabi9JC9aqtONqELyQLFZRx0NNl//4BmY8V7WxbT11CKOonF2KAoGDYZvA2CxwiQNQEcxefetI1I
bhdRbQ4/1sqI8ivU3+/6NprlBQQAwH1X2vXmosr6CitaeExkfQNu9M5yVfj0MYyYvK3hxrDyG2/Y
C+eruSRh0JCrpFU596SNOER34SLjz8gCSNl0nChmGRBzmK+jgY+OrbWzH/ogV+TyCOU8yDBQk9bl
wDCs/0eSiTbtWMW6KFzaHL8a3tq6VbqHkp8vNVz6VVvbkdI3cXgP07ZR1chv8Fh9OCaztgHzCqiH
CFfyw4Wm/tgHaR56C3Mg17lEZi6VXAAvvc0d75G1LJdMjrpzpeSLGpaymruWWzQjuGEhjuQS1OtD
MoyQPDY+zrT8RD5kJduWL5ZHpJFbpewsMIuKebOHIEifwNg8FKtNU7bBul8NvS3dzqKqoAjEun72
lfu7GyI2IzXC35qkzri8o7+XsV1PZS3hGHt/tWTdnaiXvSeqsbsWVtkcheY1AsseQ6Z4xMp2q85b
aEDG6NT0SUfu/nnudZlQa0fVJ7Ln97vt24hIwR7buEmyJI4beWTFSwxrk6uL/RCcnHuMpUtkRTss
XaPvATl9r3no18OWXp8hXvaDG2ErsLLXfGoUV38DRJl/ywf79hC0l8Q+nwgMlu9WtkwWrHPbP3Zk
TKDsTDBnuuaIci9tacOLsmDVmyhVJ3eS7Ga0+FD0HhnrBzLGfZD5kQpBoQRh52dJy2rg0NjFMWFx
zHGj6yryhlLifU6fck0VPs/LVFrEqZNb+WEXEkajfTkEQKgGKQ/L4BpLwbm/JZYhBhvKmjUImHV4
9u6WlVKgzE57ToWPHN4t1YTiZkMk/A/XY/45WMs7eEDUPAFaGSqcrf5z90fTfexIAxniO9V6Gcmr
LebyR4p0K0ENNhyniDHT4QgbR8AW/Zkb82tUe6LPT0khQDnU4WTvwFU7nJQwAAZRqaPg4/ALTTCk
IpTIjPYESbm8SYcYLnwzGRvvajPOfx5rF3SX80BNNvsPAyu4tk9ymUd+dQC6UpLXiK5OQpMlK0du
PCdbSf+8q0+DjuzfGgcLvloAsjwW2xtLdfidx6eOQnuaEsbtefUNMWDcHP72BvnjOWyXbAzCQltl
uDFEEn/xVkYSjJo1BS26j7ov+MLN8Pfa59Nzl2ILEgMszuPtotpbrL5pc/Cv6QZ2lNQzXtn+tiWU
ssz70RTF5vH8w3wB8R6aq1F7JoAODY0qOX4dqCIab7h3I9kA6Th3pb8iUC9Gal95VChE0LKiUN0W
eyNbrIQMRxfwT4KHEZqMKzn4PMDCF7vsU1PSjRiidauFML4db4TCXl1NJUwk7SV6C/LrUJ1bjJkP
cL03fqJMi9zuHgoJlvOAPXaTBtK3QhrtS/RyqshUOyJlUOgR3+JR/NGG5FznB7SFt6Jar9mGHx3Y
Ki7vcKe4KyjYwc3HDQhDfbEUGfnml6LlrIPKxw4nrnYd3E+M1n3QODfGQLrOI06rhUqgxiEVqidN
K4f0Y8PsB2zOSbqgsEBq9m4tBliVHrbCdO+n6ZJ6U1ntKIKK/SqgupHu4TagHrzJcaR0rl5/cUtW
n3ueR3B64Lre4X43z3Olg3B7jruUom1TBcfjtG1wiC9I52U13mnBPZxQYTisXcxfJqX6VfJeyWQm
LBoEy52IsFniS+YWlzPhlv1r88o8dPWxvAM1BEFsu/bcEV0sZf/BvRewGPwu7VGrjSO62zt1JQmI
7OIPgMdqrkFLMFIzRaDzlA2b92Cg6CyBH6cI+EuJpcn2woNuP6ZSSu9CmQaexkQVHcdnXBu1Ji4n
PgzvFo6C/1s3GUj80k1Bk+mlVr3Ibd77lOdx1gud36avHdTPDjL2pEPnJih15EQchzhu4tRgT7f+
WD8Vtq3ES92fL7ht974GBdjkOAANCzwXeNUwYBHy+i/tTAZS+X7p2El2LFrJYHu1bvZuORT6+Zc5
5avQ9EUFaQ/EDsic/dTwzd79km6AgRXBcW8O2NKN2+YDQ/MfGnrVDxWYn3ZznWkI7nMdyTyaikvu
ruqdoVgdlrQ3LmqU6vkGYE7UBmhuv8Sr1cwAtgQAPoa2RMaM7m6kRCB1Up1Eo93gGC6vs7zLUqo2
RJlzAaLgeiRsdQQeS4X38v0L/nNyqf2GtTdpbK0BD1C1EEXCdsEgNNNVhzJirk5yTVAWemc/GyoI
I4GAiY21WssQQsbrP9AXWuClFfJQU3FHQc6eqGcoGm8nMksHh3Efke/A7nFekLRdflH7L0BFZ54S
Smrpp3UtP6RCFGZXlW7F2cunzUIXDyFX260DIQ3rCFf5jZkrB9jOtDAA2pNIdBpTujLRGVn67AO9
6GbjQaq35DdpfInO931Uw1I8SbS5aT3gS/YHD7k7ncxUfErpLTm3U6qKoCZHKvRz+WlyQnW/cNJ8
LePZylcnRbONTSZZ6PuxzY+YmUajUQN4bFcY1tHH2wi6EPbMA8bvP1aee/bXyOGUb6jaNysGN5k3
sDG5e4U0VpCxDuZKdCWLrttWRJsRPaWJGrxTb6FnwOIK2wVFNKqzCPiKnQoGMtP27NmL52d06TmC
j81JW7oTLfy2mhZkqFZ3iMqHKqrbQSu0NU9u18QrfIBVJsl/lP+MAqAiF5k6RUA9kW2thvqfS6mS
S7iG1yjrVxRs0x7R4WWott3lFa9TfosL2jxQ6V2m5Ngr2ju59y8St4hJLo9lX8lNIKWtvqSqt3l1
WopnbFB27RJNe5IVoEnbbMsrQRVk5AEJC2FU9jevfP2aoLeWiuHzd4gEqqM9139FE0Be+WA3bqSq
FCipG6EHjCP10PLiabg0/T/XajIrKEiM6lWMSWpTlL8yq3tXlyWUKN5jSJ0NCHaiy6uZ2Z+JLtOz
WrNCSM2K/gfD5Y120Pm5QGB1lPXxu6sKKvYD0h0jnKRnVw5fRKy+0IxYb9pYLly2BW1K1Z6Z4Hxd
lLwVyunkoAGoP8aVs4KI9eL+GC6uTkTKil2td1LwVU0Uv5Lv2Vf2WAS0jipIx4FAD4+PwuNwbBV2
VvIVnx2DIxrAVePDYnvVYRp+yF4kNS9LZbYXRq7OCAL26jr0WFE3ixzUSw+QgTKjEgpM4f9PwfZB
jwLXH0nFxKVxGLU3F3CE+iX7WPt8UjQ91fb8Sul0nkw9LdZhJbx262w+VahflifIGtsNyf2Y3llb
j01Wen16gq92f7aGXUFPgpuPHUmKhlaZmwARVp5N8KjEX0wlwvIJVhyxb77HQcnhffwHEav7bjS6
VRZr5QWpkL8jnMI4Z7HvTlyO30hx/JKsHj61su3J8tDG1+4xfunLrxa2/+tPGO3nxhGA8mNJjC7s
SPqkrljc5lMFATSR3UyJNm1KP9cpxnnJ41z3bKCC3uGZAr74tojRCpwuGbjpv5zN58fYmFI1JwHb
bn1HVe8duhipXAIPOPNVG0brkroRbdzCj/IAoVvDywjstzLCLzsRj7BzhqFp//pXxi82zwBcPeCX
OG2eblr4c4/Q9bpd08gPzW0/UuR0lnnBmaIG1oL/kT0P3r3f6IM3rPyP3+PhMPkRkEpx/nmkFNnr
B9kDu9aYiHW+ilGoa23ozMxi+m5alZ+i1Nn9Qux4qCrBAvKus9gEuW+YmJ8dzvLm82QkaGe8pCTb
hMAQ3aBSsCET2JSI/Dg2OCsznkqpvPjVk1V0AAXUxO7h5lPgsM97Y4DRAo1qVv2K5V+KTpV+Rc0K
2jOSbU4KcnLn07EvprP0Z+nF/PRzibcjHm3zceGVLSBOyQEa+g/f8QjCQxN6xEQlpzPbogUHt9iU
n8JaAiPSNrG8pWR4xdRMCIqtUUuilIuHeVGMWtZmk7Elh0OS2OG59OPmvwKCz+PGgPAID/Dltsye
7VHKFahrd2GtXu7DjOgvWUgLvESHWGrVsZqc9EohohSieE/h7A1+o4YV0sdrFoyMSAwpUhsURw9K
vS48zDdWuRxy3iUeI3LmphNCnq6fBZKuWNpxkh3CjNOqB+l06wgQiG9F/3J4cDY+hkNXxMoeDce3
Ph1NpdXph5+I06YTMZnRIlla5kcqGlfueaObEopGaudTnsWN84EJzQTSnU7nbV2PpkdEAbgiqCx7
vf1Id2NPMhC6NPVsjF3AeWI+tWiMdLhpdMAGE/2f/3/PNxwLXmtkCSytHsY8f+UUi7Bvip8yRhXM
0O/eFNsbFERgE2hZXUJZnEmc1D84417crm2OJOj4dYBXby5U34Y8tjy3PaD6kbN4+XDeOVCb5mdR
L/oX9Qd6U2UMWcubuDunMUYMM8uyjuZgWQQvQeklBraCWfi5bpv06CIJKw71sJMg4k3O1+iEFIQg
F8+YWiBDibL+Tg2LpaSVBS4ZK2/cDL0rOdTQF8EgPFKhZpLlBzzhj2SgsP6+vTlV5PHRPxD5w/TT
hrDl0oT1O+7gcWiuMsq8Q9su/2+AstaZtuickTVIdS+Bl11J+WJemFlSqAzzr26CObM8yrHuojqz
TvSxiSVOi6KcG2I5+zAKJmlutKqDCC4CFmh1jGM4QhrsCfcgfRxaPnzjIbWItsT26lr68oWCDy8U
SGjW4J4BfcaRM2BfQKkxU9T031iTUqIyYBrpkhgii5Dvf0DIjYfbW3T9I/JiLycS6gBJAKnP5vPU
Yh6Wo3xN5up7e1FFMhLgi/49UpSLKQvRP0fbPgfV6jXJUjQS0DOt+Y2mrnnAH5lQaET6Obu5/vCw
k6FYCmuBcdHOWrfdlCce1HJ38Qits4l/gKj1RA5r/taORp0mzUFgLVp6BLbw/fc65N/mcBDPrPX3
Bnj8TTG+CCBIQc3XPwGaHCMGlLCy5Z6OOE/eMPdOlhLPrBhIAz7hQDEMSUIAKL1wthnqusR60d5G
CaDzeNB59nP4FJyp3vtVv8GwNidv6pw310aT9oPNB4RgOsuGXI5LxiDGKtu4mvVkvUe2snGzvoxv
UmkCuFMjrZKIugA7TBQQuzmQHkBQ6JvSnRTf65d9XWNAG3lyDTx31/xIx2q39/z1dUFBw3weVv23
sx1GvPpF1CFVn5stLu2Ybz2WwlsbAdNabZEltokytYnqpZQSLn7dM1E1BN2YaYI5vkGYdFOxD5xI
PNBzdGm3PA88wWP9QnniCSRyypd+4vYux3lNISP30+2YdmWoAnsoqy9HDDRGZvfVuJ4A/v5Q7df/
NZ8ZuFFsebIrZQswvhFfwIlmmCxD7pWa2eUrvMZ67IakCkcGHXiITSIhKw9cCdten/R/Hv9DZFlo
A1H4b8e1QwSkfZDUADSK2H8SReKSxTZTI7hGiHa+Bsg94EgEER6ubaMBFUE/OrQxvEkXV8klapds
dAllEt5yOSB3pYmsBKfEl0R8xv+ckK5Jfz+KBLh8ZFqMeM23PeZOsJW0T0ldPiKxu/raIx/A5JMW
dYgg/5qrfUG6VHgD2ZzbXl5KJuzhdjX0vSn/OmvB8QBnjBcYQZPR+LDdKD+MRlV6cTl6ky4IndiG
VOjfgVZu5O3mvWeHUDAzpq+EQ0+TND7i2aCTTqUGCkB0docuN87bk8EdeniuPEFkWDflbxo2nWyt
tY2SYvx6FCuiO56PU+gWZ70NdtibMvUlYM7pufDX8VnpvVRvj1UTKYvfxFlJbQ+PQbzVmP4yP9JJ
bzbIktSJc6frlU/RnDvuguX09c61mFzCOJdd+RmkhZGtEwwD2nZsD6eQ+76ViaJTVfx7S0nwznMU
fnNRLdXo3odnI+oKIhzpJjvMaJRSFR9KnwbVEmhpq0zUyxLZmDNJAtUkKDjLUehIS0WHAtHb/pie
Q5qMvd5f5PLwa7q3Ixwda4WkiQeMm8n6PKfOyulaHzrx4XjJZi43kKpF/KqgAvLQ2t7CuyjsqV9N
3vXuyTl1vSDnBornAu9THXuS8wapgjeukgspacd98QHgvsobdPVs0kMOAxZ2RXhFVaIf7j3cDe1n
oLXzdDcmrYSUIh9mrpCdW97QJcCxNVEZrCGk/WYh6ihdBJYRHSYiEooRGbSV1yPeTcTlHA+QtQMk
Sx1UW7RO45i70+vCWfthvoZU9g6ROGtp/9fKT3uuOOHk6E2jJD+EKRnWMXpa2C3dk5UZ4f2Uc+6f
i3FAzZCzlTaE33N5/2V7I5ycEdkJXUVbSGbc+1jHTSH6HYZ8TyeWH7GTDN6Ep29P4/kGhnxciz/g
acMYXvoZ5RiqvWdoVCoiU9CB6BRKpIiHdmhJcFdqQ10b6zmFPrqA51fB3vgRgd7YO0G+TXm4LBYv
D5kVLpfvzcB3PQHDGZ+nczbVgWVbbVo7aF0SJaQmLZf+SZeeOAJbeqvJ317spgLGR52TiVip2hrD
IYOi9/Y4Y3CMVoZSP8Ah1ec8lBzw8zbBkga3NH140zRyWuAXGgCK4sdHHCMsKg4UGgG+yEFTAHOk
eExYcAxEX0IaOoV5PZv6F2veClqXkHJaexzL62D3J5rlIpyztj31VuueqFMyFl4hz7egelOKOnx4
sNu7XiAHErkQzsI6SX6XyBpbuIganbWhQG7qWmCsnb4uZcVNKXQ93CwbPtCfedzjKqn4C7Ypt4e9
wDF4/KYUnUsY+vIk96bDeNJwaFo7Y/8we6Gg9Q52q+hI9JbkGHjl6/M41ywbsvIrAbgkSDp7qYM6
UfPaq2ASCbpMGRsrL2t5zTLg9FuQhXkIG7OnBaX878PP6aObasdElA4jJP/97AQcpIDQB2SE+TIb
v/D1pFRnANOZu5ZxbR/XB0Qk03ExAM+V/TYeObQxvUahYkjrxvTTqlWyiCuH3I5Zomj5vK4tJHXA
IWpvfO3nGNi5VQ21DP4YMbO3y4P+3zOqp14OiiWtwF2BySvF3Phu34mrlsVS6Skqw6OYSjluDJQg
OI/3mxAS7pMTFiyKJBsj/GDzHmAWhlc8Q3Tn04H8peejnX0ZtAwVZsrlZWlhvPREz7LB9ZmgHXLv
/GfrqKGhU/mc79FQQwFxTXvhxq6ORPf/bguAzRFVMlmIeFDEb/NrMQxQgRXyr7ZA8T/vVB32Pjrz
tv2AQrQkSz/+Kto6c8qIi5pr5ZePzALNUmEqQ5ojhpCXv8jPz4a32uC/N79ov+KkdulwVSVKP7U+
26MyhnFYrNhKcm7OJxTFj/TxducHcKUU3UczrGxKftsER0oHwYd7gnYP6PgCdIkKkf6Q9Na7lHCl
vA9ozp0Q9vgLe0PkazsPQO86HNNwP5R6n3se/pNMWwnO9xdQSZqgeXnkpvdOS9RLyTUr657KyHta
Uq/y0NBFrG5AU+qQfdBcFd+itpwuQMnsGYRFD+18oqKKO5NdqYvj1yRor98HmGZr2gZ9YmGHC0e8
LW2vVi0hNdHI/E+xmMkLs4043JdJRgTTfMUBppWSpkjEr/vBH3vbpsnL9BVheoTUFrK0Xkpo6IB2
YUsyZW8/OrSDOgvMA5Zyw6t6pr2HhoUdpioDCp6Bf4bWCYfMbH/Mk0D3AuhFB5GMTcRBLDHp+cWb
7c/l2imeGmzC8Qc35MQkiHvsVH2rXXwUqmg4drR+XHkZRBrNVKoV0aFCx6WYQeQ4m/B+Tm1XI+wy
O41uiOwEdBlZiG1wcRPnDT68sutKA6vaEJd1EJg8sZql97L2aUQx4RyeJtqpp7hcDa9dmCOOVF0A
3iEE4WZ1OqWHgqAbvWZrZLz1JJAPjgIpVP3EBKgZqySvNJ0D/03h0kCE2PPUQ4X1X9pUk79+tW7T
mtsUwh5Q361apMGoxQ0p282VJZl75gynOkMwEQv7Lb1pY1rAjs+eZuWyLYmPBW0UxwJT10mRqtOo
bAu7lzUV+KaVdkyOPaq7gqCJo6Fm6vcsfdANwDIWmrB2cWDT8p2RVphvR/mMqy2M5CCk3euVZODB
oeGZLkHhJSIl4hYgcuBa6KzFFGcPlgRsRx/QkQJQZcz8eJP0hYEKXvifI1X+NWjE1BVxvxj7wDk6
/UqztWztcGmFYg6WUEUwJZd+PKGATpbI62jA4KCGgbXUAY9iPrn31Wb+4Jk7g29LVPu7TIH6kOaR
EmGzcsahSEfBTptPW3/Oizx1NQA+a+Y1fK9N9yCh4m6ziqwd5ct05KkdzsZPLYa1uuLMQ6XPhU6X
Fzo2nkBNln2Ml3Yvx0NFMHm5qGe2CG+PSG40vQgh2vqtfXfuJQxRWpmKXfwVUBTnf2MkbkJSM8BC
GGJTaayeAqqOJXyB1MD1O+A2NxQ2YIs1grrnC/jRiCYQpRyWtsy/OZUwoWtXnZOOKLQ3/xrMesNI
y7eTYThk+IJYLk/g74/Eu5dhjukMi2SsQjXjOyiO6Tt5yEpeEqnYSgcSdAeNyuxcifURuIDuDSgE
YjoWhXJ1NseYkDJ0fyf5Qq/M6zP4ZjD0UuQI6FVjuYiCqwdCns7wazZ8QJ8k16FkSjLFyvfC1n+D
PV8McAIJ1Q8r+qzkao/ennegjyHusg9e5a+n/4LQfIlgxKt5hTgcgirw8X51xNXx5sfmuC2rLwCi
0gvC4iANVt5oNuPlLy0VPVl3iFJC4m6xUxpbGVGKfldHWBzRfEzkO7g3tE7qSHXNSzm8r12PQjQu
4tXU5ueWpTknLQsI+0bJ/lZrurFSibblyWbhg52ltIe7BouhTSLXIhD+6cLckmPDeoXzFbTK2yHq
/EiXMbicPDB8NT9GdqjxzafRkjXhY038nPbo36b7cptYKkWffDEbkHYV6gJPr+KvYBQb1K8ZDUQt
am6xsm0v2kCmzc3nv+DBA0zSPl0Ja1G0ugk2CNxS+dS/GkVcrVmZoXVGB5FDgyZrizxMnPX1uFNz
gRh6nMNac4rq3MMp/m/g841w5tdFOgdrOFTbbPujn9jLTumLghgTwkzdXE0Ub6pp80Fhk4M3/j2I
RLeXM0F10ex9oHECQVPt3vtuLGqpFTwNZbqHdoqspXpZHIqzn2eCtYCko8/Bh5S4QJ7b009fqUe9
e648PMimeMeP4rVP8ak3k2pgHfaBOvnzCWRpkuAsQoDS/dNw685th1/kwXtORCZUDlJKhhg4Fo4F
izIDzj/gr1WzqNbQEhQsS2sdg5YSFCkvobYl6KDHsBrVX/OEG4uLUDMXYT6FAeLNQHTiFiiInOIQ
awnUVWcIQtX1+qp4qf37U9FQgh5kpI4gdAYOaqzaw+VBysHlmVImXalGgCJMYQHrvu43WXWTNki1
+6l8wdK0hqd96B7NBJgc2vG6UPXibBft+QEHDAF0Nq/Ny7Y0DJiJ/YqhnpYgEiJK4rXGobzup3Q+
nVgERa75qMOcufIPvFIHlpadbBAe0TcOlPaPQzKzPIYEfgtN7Ai/U/EDvWX8NJXLPhS1oeNiMURx
aqghuXpU6UX4jxLt34vdDD4UnmkI1f3OppTxaVIX7e6nHO6GVzaF7WlOF/BvRiGVnLNzDq/90kn1
K/zgIdxaXgVBKXuvm8zA3n+MoG995yzMBEeglzg3MpgJnNr3a3JYFocMsOsnTCZxZw6Q0K59EVZO
O64glWyn4r6/IEPzCu0Gwe/GXVEIE4OevVUFFa4ZiYIbD/dFyIF+WwNZlQORC8WEBzVXT92BNV3O
BqyPmdTgH/m9vJdJoh3ewzV07XgmQAHy6ssZyQUd5NmPZZ0k3bfL+6OuDskHBD2jsterDl3MtPh3
N2e/8GgsqdbW2vzBmKgUi8bKZN/dKadF7V16ZZ2HYIcIboLE4lmTVM52z9nZGLqjoaH0gH1Lel7Z
nYEwmV5nbb+afp2DKqeoqgBUUigh+oFUn1zHfFaxlWHwK4c6L3G5zBR2rabWxZIdGp0oVFcEI6op
YEZ+pcgUqsmtVN0I743CAloToSMnxHdCbWlu5gcMi3GejcDQtkBmxeDbtS6JkAJ/DAUYaAaxsJ4l
j0CcHL/DZWU6DDAy0hM0P+PFuRnc7KqKDW6jsm9ftX6dhRjwTDDnpXoJHSoyhdUrLuqgF+a+DbDV
7iagrIMS0j16/Vo8szBgqll9RpPh1fPzQbwbODezAiCPutwkk55a2vOBx2cpdxItGLkGO1U7BxkB
2HodaM20pdiDBA7YNhSkbtTXoebbyLADASpaFs1XDWluQHHiddqnXhypkoZRJvXSa//V+wLQvvMm
YqcpxHQBZcj7h7ulhr+YEt8ZOLVuaVdX+9jKo7AzVRmm40MF/DGk3xFrynLAyvtT+VNGJphCEFhX
5DSw8F1CEYc6i9x9W5lKkY5Z7TcLyVY5qyOZcE7yIxLL+8g6u5795WfrWV8SEknPtC5mwmtT1wZw
7R7xy/wDVH26D0ynbx3s9twhbfdh7PHuh+SWwC/2itTLXVi4AeVEIz16AA/sbWEnKEy7At5duJQS
eUk7NjIirWg4RRIt+Tv+JskSVSNL1p7kU+Ef1OcGH7qKetSXaIdxaH9FcqIH/0qczUHGzBlp5miR
8iPZ9vuzR6R5o1Sl70qdpXb82ApIZTJHP2Gr9SupjvlBj8hFYLFWzhxcThm0zO5XEt7LSTV5jQbD
xQKpxy0dFMPAkxHagexLVVENIoNkegpIMoR9JqVAYTZy0K6diBg9l7pO17CynI1hfOE1tXWYEnfa
gwfwvgLsc8IDR+FSjUTp2GpDOGDVjFtOQ20Yz6drBgfaPVe5PSpVTcpGU5L2dMx7lWFxbsK0KZLb
twP3FSxBE99HtKI8lI/tsKhkt3Sadx8uK3DcRqpCJnpZDh9XIV5JDpIg+WpJnijzID0l1yFNRCXR
jH3Qbs3KmSqyGJyGvWP/yvg5j6UJWbJd2MDUzmeesGJ+RAmREKCwlXnq1GHCywD4husHdBzfQ3uc
ZZlo64xg84R+RC7mREbw+zD9GyvmEIXP5ZS5dew8fAXJ0cDw8SnYStQ30gAv/OSuYfeNhKe0Xy4+
QEWoVOugJ9r6i2EmMKdpwEiMY7CL5OrWNZTSezzhZjZVEnqPWL2sgfxWtyn62S7ir/Wb5ZWYc/Gg
YdyuthCfDfze6wNjsX5Or+/LWoSs5W8g9tdGoAZ3mq5Q2hSWEiDhJbsjicjacDnLxYHhscBfkWCs
eCB85B62yr3NUvUhJ9DFRt4jJyQ7X7U5USDs7h5u7A5wFPEigtXkUfvBdZQAQp6UaHeS2q4jC+Es
g4nxJMd1LF0mjxknL6TjicEmf8Bfl+GecMzgsq/3x9U3Qe0D4J1jIPSCZ9CpfXNIyJ2xJYExJH/3
WtIBKnV+tbhBo/Njx8W8NSogGFUZER6Zv5j8WLKhtDa82hl3TgdiTKf8u1eh+ugJEWk1HGnA5JsD
adhPfbp24dcTDEJUSLGfNUCsQ9yi12DiphwyvRYvwPasf7TcEcJlfAk8dUbh/wZfEZAnplujwvoj
oRSh45UKW35+zAtJPx9ULP1bpMf7EUO5mUcfDrz7OT7/l0B+xWqAvOFxRgauSvntHmCtHGVw886i
MqfyiFyb06lPAD6hQ0Jz+5mDVP5zydBu2moulkXob1j+FY0lt0UVais8zo1oLfMQuNEAGFdVmzKL
rX3WRZ8qOs+InCumaDJN2oxRYno0H9PTdT1Rlu82RZgnO3HxZiD+brpzmyJVfH2kTE0QomYw3DFG
N7TwjZ+zHlp4MFKVsNIT7jUMQAIpKfec0A0HJZoKAO1p9W08pvzyjV+HUA1G6AD/Hm/ZrbZ1pm9O
15LuWLim8MI8031rmMol2u6fp/XkfWBzEh0PiMP9ttqJmlMFa+m2wp3h6FUXmIg2Bz2/BMS7h1in
17/wAtp5sV/e76ODqE2ZavvVHIHqwlHK8db1f4lwdEaJ6+aVUxQ4cT2SvwtL0AWYK+UCFIH4fRGq
hFE4HyzIOodbSiPwm50B4zUUKoPITN5/Wv7o7LXRNkPR0cR8JVfNee2cX7qZaarqdLyjl4gnfamj
VLU9MRVY40CvKo7RBFQqZUvSoWqJHzu3sSoFnSfdQ9DYwev73Up+9Yn3Lim0uCv3GbdKTl5Xmrhu
3fsmaP6PXCdezVj2rVkYSpgfC+sMF4eoDpkrbFlxHZDKJT/lfg5HfTl8EKks9CrtdsfHMzY2F9nN
w+J+THeZ60eNXbxJ5Zs7AlPN5Rvuxc61uxt8xFuvACR18yps721C+k9IzrtTiCx26zdfdkV6gFqM
MHAagmUQqKNGOl+P/qX5z/opL4bAVp6T+tDNMDzLiEZpTyWeO70C//gTUBcXejPJJ/7graJdvKif
PC4DpsL5R23pbdMPHnkcd+NfViLXEf63OIf/2Py9AsJfRR4VkobJBxkOCE5M1pm4beyC0AdzJ4VF
nkSlLfUU5c9J9QJ1+z4paca3EFignQ3W8POiH8Q+J54b+Hi7xj1WgqP3lWLBUvfijymDMjVhTmEz
7++z7Gohiw7CLFl2z3Ld3qYmBO13vJFE9erQD4bYBiJdtsPYcADTSxIr+QdM/AD9TYvBRXRqin8r
N8SAFDGwBVm9er6fdROAkWdWoP4cuANL7tvjqRtd/i22MYiZTvIzhj0JKUYzdb51I+Hi1Xm17YO4
mD9XYgwWW9HLVOqduVXWYjJ2WwA1mAvnGBoH6kW7xGJpkxj6vtZLT0wT/81ouOR0ULZIuG9KJbcB
i8kZ8jytX6CCH1lWy34R9k9LU7FauX/SX5SBYnR6a+89POvfz8KZZWv4PRVC9VJBdYB00wwwFzKy
HN0HsrbYUL/jDrAXDHstCBo6PUXGd5gw2pQNaTCVIL/1jeaDwRw+PK3nTFjLLpU+Zs/jy9O3oDma
OAQd2UCDw6E1iQczwG66ofNHKLxhMEgm7wpoPhBmcVHI/8fMk0ZsNB44Jieip4rxgePe/PY9UpOb
oV5yGgPVId5mJKIaPgrpGfB1GWS0Bl784f8tgCcyeaYTgNTkuQFiKq1UAMNmGfusg/JwnZgjcw+s
qgELzFMozTvGi7BL92fG9P7r0pdozLBfEzMkf8NdKEcEZmGnIcghONYwt35gc/jPD0W5m8TKxX2X
eHNa39FMSPFA+8VQ1EpLx0omAYgAIKiQn+cUiuGMgtYKqBmN2zXWjMDeW+wjXX6SBJhqrl8saFW9
ce/+X5jyPOnKMbj6j2QK5t7uxrsQ8zyjTnaM9uuMtbPfd4Dpgqn3fhJilAJUE3La1APsXwK9/NSd
54bxrpLPtkHmfAzB+W9TNF7wyi+oj/3bAUfb3Y/uUHVHXIkNCDcTj7kvUQwFRu2CuAXrPTT3BDSH
NZcF+72bfTiHRPh8uGgJh46eccUYy/9qCsxOKSL6qyBBNiSGKRJcCRIrnG8oB024wQdGhBoAFDh9
iSW0ZvX+xVGrwE31fu1EVe6FVx8TdW5Dla7x5iYMCgUEaf8w/3vG6kcyf3p71RuySa9TBSlCxrxv
HXO1Z12brlqN0oBHayqfqw/mXwGUFvlel6bB3jZMiu3iTKdKU8KunAUB0MJfA/0n+D3WbnJrUhw3
IO9NRyystmVNP0YfcrCuhEF9l73zv4QlXwBYEGZjOScfcVQFTj0JlAme8p22/JjIRNoKkZvyysLG
wmNpmAKpaL/Nbp23EQThQ09tVt7tJ1RNCg5nJ/RluYjUx5xuE0gtY2dxkSqeNcoGPxOql+QbduBN
ZsmUUn6EqRTkoAdZHhe31CaUEPQ4zyGtH0YHHE8w8HHhKC0BkuT1uDRqqVyyB5Q1Y2rmqoT61iBW
1FfGGzbLjC72f73xQtTd7XVZSs0BjCbnz66NEUwg+IQaaBMYHp/ige76vPJZjJE/Fv1BJfLHAb62
bUBQo2a83IL8/eGNCTjKUNG9FuIKxeUuqiVrJ7XqXXfdmPcQm8gMYddxUvQUIpNUk8hOmXxkksun
fm8ZByVNKnFGeWcvaDCYKiW87HPZzyts+HFea+Su0fdCkUvyzBKGQ3TeOSj9p69BRTKmIWcwT97q
okspB1iCaVH3sKtcjGWEgBb5BBe2EGrcUjGQubfGJuuqODvUiJC33twkhSBylNjlwTHYaY3sKTUw
NyH0XB217sOuMBigRZW7qvR3/HDgD0xx2GFl/9Oq/8ZBMMO2M4VvnVCN5ZZhjXuPui15JegD45He
qaPCa9qYo7ANEDO5tJOz//kVpgz4+O8nEt1cSwWSXAphgJWIiOU6JDHbWDnyokt8vHmfIHY7C9yQ
G3s+zlfRDwV5mkU/P9FmgSiSzzcAp4Z+RaQ+/95CxMrxBaZ0PfA13m7QhDBcsPebnqUUm6bGp05Q
Tf97/vN5nFpvllc2bXIxGQ5ReG7RTdN0Bv5ycAnmAxRJIzcTHGCbWo0K9CREAoLRUxY4DURHbs/0
2qD9LtRZ3NzNrG0OwhAFAypEAqJHxqmaUA9QMDqFYqALzuUJ5tVRTGDn5TcZaz1BQ3YZl5QROU9W
+t/mFIHxmKM0x/Z6Sr/R76VFsFvD8YBVGjycIGbL6Nf/hKr74z8C0zSkpyW9d8gLLNl8NXjnAV5S
IOmG5nOLU+ljOcfTaQGIvw/j+jzrTQuGN0HZgtGfDtE43OuNp7vyahvCd+oQEGP5EOS6BLauJsDP
u2J7jPcw6iPw7MaL6k53sWSn7cZTfZKAUg8iQchr79nSkNjXSQ9m3PNjDGK0gLrJTsAjFoKVj7js
RoM1aWyDhdbkcqj1jroRRcCZ+4I+8X6mYPe2TOt1Jj4016XsyGF0KxAMMuPDOlxynf3JlxUp9tuC
n0IQyTq3D0AmdfXvnrTylfxsA4OIVl6QkSyslMvWVuV3Q7HDAvvrmprg7HwLmP0VRqKdMLiacxBN
fxQUCYnLFvJvqedLF4GfGC6On+WIBFir8fYWsrHngiq/cJqBD98nyGQ2Y4dhdPrFOTFOxdSEgwAG
/83cken42YlmskPyLF109ha2UH9KkuxsLx5zZI9VnHPFj70ovuOlo84gu3z5fbp0VGtn/xC1b3PE
dyTuNG8A0aDUhWUOVJGpRQg0doKYKDKl7wXEaI+0VZobMzUzwgEBQIl8j2K9jExf9pVVA1OrnFp0
HGl7Yd5pE5mEdXZIdsZs8ISGKDQ5NBX1GhhrzHGiTbQJmvmRNlA0Y6tORRC+1WlKcotnclZpovOY
N09f4riZmI8E8AHiBMbU8Ii15s+P6aEzBQyenBpwygc8UHkFywhksigLLCoUa6f1V4KwAlGPmM5+
FwM91xhD0t+S8J/5AUe0Pioy6WmXLU528MHOrys1GVEowl3gmGJEeYYSIA+8eq4YX14hzJGQ8ZSV
tF9Bw3gDIjQuQFegwSqCI9HvwLiwrZkX48bfNVQV+EOt/tDVvide+2pvGNfLgQWShZ4rgGVJxJmU
/SOwI7lNseGTRZi88ZQtUhITGrg4Au7EHqfIZQg2Ex21/e2sNXUpVTegDKU6tNZox8YbA78/r8Rp
I2es6+uMaBUiaPkJpiMZJODb1Ezwvb12TOzuzaMSLDwgoY8nn8MMxg59B61kLDBWcA2KcJ2Z7R7S
QTzyJZmAvxiT1nkJPylrFB/n6M6s8AhIdvWeRI+FMVimvss4hgZ0uGxkiMKi939QB4thAZS0uSM3
6voAlzTDjKv7r7hv0s/Et5YMyW3c2lQnevflGCya4AcoKHRbaVkhvwy8pKyoT2hcflNzT4GvQP5R
rnyr6R2GlbteuWXMCGo3oZwnLTEjYdC0H183SkuYq95/HebvW7G4i4h9jG68C58FhbpxcyDli1r2
Uh/TcDx3LGhA5XjZTEfs4G2GBN8TuJozdZrSa8CsWgHI/98UaJYhP9/CrqABy0q4ald/knfCqanV
qM8MZZy8dux/ldBz/9MQjp0IajIYZyEGBgtYg7R22kvuoEVRunbArJTGN9WhlnuXj2CDKRJ0LtqI
347kKlS9QsAcaoXsX2zs3Fq38xl3huTWSXVa5dhwm5bJri50jJn/hSI4U46+/10HMvDZrhZzGZ5M
Fc3PZz3247LPcracWdea+0a/Wq3zSPSvjByOSjnBHxLSRNefxS4IChDh3QdJT5e3e16IHKkHQwaX
DatmF8/imPcCalpmE33nZvWwxnUbgzZPgTluAMDuOkP9UdvGIYtIbDTzKApYOM8rtcr0Squloi7F
Nh5xFTCpT6pWdMmC9JWlaSrpAHc+N7rQdOuaFe1dODJT2WhEan4cmEqR7eAqv4gXKNYaNiFQP/0/
0QOB8C/F8m4u3FGmPE+t78cTgTRZrEIUflvZMT2uTDHDHRdR0rOv0dPdzgm65+XUmZY6WvC28fWi
UeDdBNHwGF2N60++m92T18lQ5H6tNYrIsT+LS1aVBQz+fbZXPZHaUgnkneqwE2/1GDOuZBVWjJMp
usTX+V9Vd8mXNAWsedhPRdF0LIIuImtn341A9y+ETBre8PMi23BL39K2EupKRQGh6BQe6EgN1qpS
oaAgoIykmH55s6ARCxwIydGx0WnNtLWKh3sDqK5ox3Zg8S+qPq+fjWoxpSY475GRQt8zNs8auO4k
GqTG0XYbur9oim5EjYdum8BF3Fsf7FSoIE1kLl+VUA17LRCIPjZCUYDOwSgj0soHSS64HyiMmjvk
8K1XMUNzfFE4E4g/ACqq9zaFdYYdSTYVj0+y+Rqqi5RNivatCrliJ1PvzYwHLi9RuXq9XUlBXYFM
5YxkM13jHCHqecnddwFuHms/kCx9kuG4RZN7pb6Eh7pwk7b+TCOOoiAQS0Z+aLewWNwf/zzmeM+J
Dz3Bof5cbgdzEJ+tU7Am3DgVco+hf3z1DKEy7LzBOf3NGt7GmiOxTkQ0lxvinG0XRuKgIahYbKrh
HNKVvF4bWqgBDVpCBzgqu8mHVPIwe5ZRPVN0plbG3szUa7A8QosXj0yF/vvJ1pH54jHe54m1X3WQ
x7IhDdMb9RpO8/dMzYmdSp+5JZkkoM00xKoM8S4DKVGZP9mkRTilWKLaZLyZqaIO+TQnFfSZs8lT
wsc3+s7ITwYHwmoFY4A2S3Buc4G/u9+1pcMWKJeRkpURHVmoisOl7Z7rfhL4Y0WAiPIW5GoxnvzE
KvDAo8t7hCk77VncmH9uvJUusN0+ofIJzLTmjcG8sr10sjr6LAZUTsA/+BYI9Db87fblji4IWryN
aTwNioSBQy4cMIIzYB1DlcZg3PlIbRsxPIhJkCiIjsWY0vZxfUp4yhjyN58ei5U+qO6B7td3tCGt
GOGitDVvIVGU2AyaBOe1xx7LSwszGcMago5wDx+zK/ltOh53L+3JDFOIUX5kuZ5qDwWcWoCJKUnB
bcVSQ1wOYKTk1B8i6LhFGkTv5ICeUENAixCs8BiQjQRifhqOwgdQEgfM/p7rHd+a2xGPpSEbmVrd
FJBVI8Pg2b7t42LY/ZlpLzxxYwYOSCwqPj1A5pljNEN6GW2qtbbpEiMD03tKLr2myqU4VSw49UBi
Jx9n/Ocle0MLawg9sX31xpWAP3QAL588Fxs9wKLdDBFimJL4Mcl2s91ydD/8iMxqNnaGh3xRIDtn
uM/MArd+J/i0ZeS2KYSlHyqQYk4apFAHSWrpESOUYb8Z4vS/yYYu0RA1WYgMbU+hR8I0vm86oszZ
uJKuAGwRlRaLaDvwq70Fe76pTgbvZ6LXO9j+SnqLF3gOGHHJ6yqjrnqs7GyJ7otMhm4XS7uGtBOb
ZI0Oi/p2+W1K8SbzdoNrh25CAO2xXi69Gphhenxpk1SC4b1tMS8a+WYhz3viMucVaWQmE69Q57Bd
ijTAVgzqhOO2Ku9/MOH8l8wPo6+dp8Njo+tLJd6aS9kTI/gvY7IlI351cxUvsHDCV7gZElj2A0Tg
b3VnMECH2FdwlRhWJJAaDtuocToXn5o3E/sHmuXYaBfWm8qBKTcPGG1ydJ2sq5KBBmk7nGk1LJQB
qDQlpw27kJep/kUYl6/cBfOB5l6/66lGzEprtyZk79Sd57bVmgqwOo1U9mLX1FJf9SOi9kXmLpWj
Twdlw7XkVFbEyx5s6rnIfSzGxsxdbwXfTwUw89Gw45kxU8AX+OxtVqsnh/z8ukzZ4yAAkkzQeVbE
8aMIqFQpPczEkwajnV1mYBlK2IN3AfFs2fEP5UXaoOXSedjhVfj8JF3X7Ju4h4rX2YndhfdXdOJ4
HgwGNC0x7Mrix67tIRc7NVIWE3OJ6gChv6i4UfoMhnacGMXlKzoRSyOjtzvYRDuGt3gWIlI9SACo
OI6kPeMx2H5yFO4yd9BW0vB3pPyTqu6jxs9U/aT6vOFslJn/DFfkjt3BTNDx8dXNjvlGnYgF2W3g
bbbdRSfXL8aabXzVM3VzCuG+k5EnFTx1WXK5gpqDw6APAS2ZHg/NHnxoysDstGYtsUlJU+knMu9S
Tdqa8N0Wv0GlnrJnbqrBDUGBKOM36rGuw+OKUYbWiWqkCq6e1wmwMwUkaLqZb2vbeKp+8/87F6A6
XYMQmIiU7x/UuIKq9jURhwvM7g2DSLkxdrL7OQbjrtFnO2eDHXRd+6u+j+2FBv2xs23pMeMnxwGm
yKzLHYM/uiinG9oX7sT3Bfg6US0r4Q3Q3xRl4EEYoELshei/6IhlXRAoXCM7Xn+XpAg83PGgq/0B
pv8O6ktAIVfi08vsIO2xyXBfCKL1PDJYI67BrwNVOazkwJuUinrHqDcdANbVs1xtbXdQRnvF14+N
P9A5/SgASCNtNpw2rpEGT4lChV7fWJt6tUZ4lD7kQ1KxwT/m/uDR4hJVkrzcLpHX61OBPfWPfLhB
lDpLOlCyK/oxVDiTrs3SCXBFSysgn6uBSae3I1/rKjH6ENg3dWrMdsa1LLdMafSeufLLCsUICFmj
lzo/G6AMHhCTNkc7GIk4+pYye8jV9Mri7hw95TKQkObeQS1NwrXkuTRlW1Xp5a+MnQ2IEpQuiOtR
pWFMbyYlc0WYHj8rVuRyXjMEKIid9wxPgFi/U9YN6bbjX1N5un+tWmLzxl81xiTipN+e0Z5VU6Lj
qSCAGT5E4FfCywRGfCfs3veH/kQGoZ4QMu11vwEEDbz+Fq3qlFZ+Mu3t12aH55rZ8mMiJb54IdLH
vTH2DxnqYvNoI+Nxo++y5++72KK+a5iT2DimnAFCxa3NExkoJ1mXl4XkSqStRBNDScG6zQ/maCFi
69fPNOlBT7rF43n0fI7uBZ/AWByJW/ljoiup7aRfA7EXnKOkh6j2mDdpRtZSQYhAYNo5ZmIRW0Me
ha0usKo8iOnNDrAfl0zwoVXUbyNRoBSTd+QS9vue2JOtveyUE1S49qiUyDeDoEjxsn2/WEJsGlCi
pBLqwgFKhpVa9qPiK3lk1wGmc5b2kUc1H9QfLLDu5x9rGyQh3E0A09TXgQn1N0k+zXCAcf6BjKyz
uQ0nvupjYwR4/08IpabstTqAJDxWNWIF2IfHhuFC5WQL60TSanrr4fw8hUtNgzYG1KP1ZsOIA+vK
MbzTyxrZ2chItrumr1r3qjm45GvLRDqdxxpIDjXdyaZn6EBCAbAUKFW2rkgKXEOjMfvWrUXFRiob
5r48mwXUQuiTM8OQa5spnTwZXb4S1/XV/uiX9OvEfVXxpzByLSAis51l37qQFXBaoUAqZOvCZ/rp
lOXQB1o7SkS1O3cxnLdzSqQP4a5KvhHNQI/ktaeMpbrZPZDJyyi0pp9fIXT2tEtNZuRKm5ilKliq
NibK+8r18doNOScdltl3bW43yj+gyzsu6NoXkwLSB8UjzmJzU04yCeNgljZsKaAvoPWGfHYwR/91
uUc9PdqYRAIA3fHHyZgIYLaHx+h2d/kDz7VO18dHJ58BC48/gble1acriI4JIQqhE+TsGq4noPJY
907GNmcGY8SNsH3uzufp9AoYrvjVp3T8DWYZO2jmkin+jHX17MkPMDLmFTrKwiKDm0PEsKclNJ9A
8CAJrRjuw16e5NS7MuKUm+4mxCmqi2AlpCL+sCJpe+WGQNIsG92YS9+1avTjzkrd9r4m3A4h9dNG
y0T4LLaz+9N/iSj/yQkFA4NEYbyUH1hcBxVG0gS9TSBJmC5l4ChhJjlfHLKyyK9X5Y4iZbfD02yY
cvFMHJ1PTlYtP0Ym8OJ0hx0A7hO2idF9xajGzfYQOAZOC6L1XSeoMO6JmqqvHN2S2iNDWNlSGb2o
6j3kexGENfuSPiF32SpWOD2ylHw+7NyjDr+9bdGDWGi21lU+aFAxo2aY1dcw3bHVIsRl1ltl5ixM
uFUX8xQQrreDhpQ++c/Wwvtc0m60zufSxkrdQRmuyRmuPlM21fLEHwXm0KceEuOuYp1acHuuUuZr
fUf01hUtMmGcCZTeIioT6XEajVeqLg4GMuUiM6INDlMowp7b2PwyFYUe0Sh+C/ORGcOW5RKu1HF0
TvRfcid5houTo8FqxDgcj1xMeRYMPdgJJrLnEHmK+ciw8ARzYuhbUtkjQf/wKFCsAtE3hFvYZ7u+
IqczS+v752ymfHn6+ANXRYAjk57RqHVn0rJ1MxHFYzAmY2nQESd1hzw9ts0/hk+NcsuwbAdcANlE
Z85hERPR3O3rYq+QMn41IwmUYyPNDMwGJ+QuJSlWoBrRanUX5UeSt48+lDzDTm2xMyP0pMNl9R6+
TaGIBMAhebEFexVwv021Ad0SM9BCEypJMN7WbnOxIXhf4Nt/Tld2rfOV5ALiVrSF1OB53n9jOn5j
WtBhekhsw4dl0Obxo7TKCrD1TV8w9vCIHfNmyLnIIa3CP62zBtxUFGeUzkbRYlb7+K7epnIXtKdJ
tpqy2D3ZJBkxW1RlzyoytUDIBlqYLLke5JUJsws8m0LgfRtAU1UL8txiXMQf+zoXIIMziBaUtVTg
MXo64HOrjqgz4IApEdeA950WJUnm9NwIplW8G3mfV1b5f+l+xq+9MSYRBzws0MMa7QRd/s2ECCUb
D6MWbt3TU1cWBSXOgzAlgdXSlZUzURBHIomz0z30rUuU2l3UI1wipoVLYsvKHQVPiMuDPUDK5gfE
cDdb7YCtzgM9VxR3QnOGw9WKuCoeRdWiuvwOch/vICU705U6VpdfFnNvkJbzfKdqihUN8BmrqrKp
k5K2sJ8iFD4COUu3T2sJyYvwMjQhJqBHcAwaN9MudMC2fDie9QGe8lB5yaG4rFtujDsl6VUY1ka2
0eLMHQksd0u9BvilsV7tVpm9CgquUKlkci29HkdtpNmEggiiQu4cHSIAmnQ23HWKFTpRpuev+4YI
TiAJvcTdd3WkwcGj9LJtxC49bjZEySjD7PBUlhPrvn3dojR0WPvP5Nh398run5E4mTzdUqax1z60
BLmALS2FSIsvBvSmU8/6K8X0x5tDc0M1A9eASPGddTun7ekFEC1GPqrHkgqaFQyaoF1jFxlzlPtg
b0KtIoNyr5YEof0Jz13vnBMmz/z9DWptQEnrQaakDTwhPDu5ytKdTs6r2RYLSTF8/XvNEMOoXe0O
Hgbe7Ke/ZaCJP3xMvVU2LN7d/7MWaMrYQNf67v5/t4ZokMKEs/99Ozlz4Vs0o440I3EBU1zO6KmI
UrasidGIIp0keQra5L9Q/7KgeU/UJQC3qHWeVu3XaYOIRj6ZJ5O2ZqXeCCI9HdMbXQj54hBvfpUN
su0n+dXesreH4yiM6zR+N2iMmLkvBK3ATLq0qQFUnvAXPnGaaPsVPvsJXyPuEtCaJ690mkp/YQHT
VufEqGPzKonOr/lw6Pd0GkTxUpv8JYwrWYQrv5zdFGX5UXguG7n3shL+ej+sMIPkvD/jv0xGgtIJ
Bk5rgbLgV7IupeX4biRRXUwCeBnjHl4DKv+CG1AziewFLDJ+py1JMuHWU/bbH/q9NBhotF2RN3ib
STCzlJIRcvHMj1cPm9dPMHUOrX32pLIA8Q9t01HaSne4MToOvSATkJSovc9vNQWKpDYeftYBPJYc
kO05nrKgLI3bjoZHpcW26HcawXi0oExh5jl+pwwr11A4w5eusoC8wbuFLX1smz3hlzdXQZ4tpPtv
4wgKmibknvX7sFVjjmSBfL3M8CZ+QRX90KDI25Ld/Fpw1mfCZCfB+95o0snYRqRRLFgXK1pucjhX
oAFgJEiXHbFLXYE2ucdFBI4N+sNICvcRrUYG1nAmEK5drtV1e7eHs+daECIEKnDzOYZ0CKNv7Z13
Mfn3DjW93nDPhFPhetyLN9vZ46hc4JlwlQPr99COHdhvu59GpTMOEzI/i3GNFAsjcI2/O/6x+LPh
OYLbMYFF2kc19GDDgpYhRf60EzDcLyNNqHiKR8EXv9NO3u56knHFwgrh3n79sysCuMO3QOlXxNAz
Qu1FVl/VZXgUT9dqbUaj34+RxXQaf4L19H1qsiDNPQK6TfmNYVPx58KHPLjL/eqLRNjuFbPBTwA3
SZklpJRspfHqhH1K9bN5lRBlLNTcn7jRHcuXgN18hUk4at816EQDEfvRdGPn6bkF6KQg8mYkPkM+
CWLbXltNwMz0k8T84AdBg7DX39kjawVTGcb8VNw4LDrz1+rAWC6fd58o16L7oB0o4QFNqtSdpuEN
365B16hqDQ8yrXKWnS86TO5RMenvoAAiTTeWM8x5LYguEBXiwtprfbBZ4wC0jqHd9Y+1AFgSmF5k
LBLSmp7CLdKVE9WQWlRngMUHA0wLM5xMDKcouZDXlQ5Q4CjS/I03rpiY8J1MK0hxhXhGWauca3Vf
Q9hZ3jRbCWXE+b8X1UQxHMWZlCAx5NM/w0I56gWr8CKHKHHKsbOaytZSjEnDXq8xAnCONS+BZ4Iu
o4phwLfq7hK3GUDIje/ICcfWFmHnAVkjjT0Q+5yadcG/Jud1df4+sNqfSqxyvb+84hsGd5lHDgDQ
Lf3mtg7iXb7TVYWLTB8pV8YZ0bnTIUutUrbKgOGu1qxo/WrhYllE3F+YzLzg04b+asSYLkrqnkLQ
C6XtgcAQBDSQ4/eQno60hDNrNcAdx27zql8jSt3U0z3tKsqzLZQ8DGQMrOlRTtjXG+8dtAR6hmf6
z7dXHMZ5sy0DK6yUVNzZUxuuGqUcr9Mr5Z341NDTwAy2py+2q9ElRAkjy1vRQGfBCLdn7DAQ7E/F
uquZnjAT8KddtG1i7LQ6d0Km5R7Sbg+oGEXLS2RxmyMcS8bis2TgLwDeQDaUrI7sINZNkgbOSqqY
4J0vs3wTiaX5Cf/BKPeHJTJ4ahhtrEdtpJey1Bt5mmdoqKOSEeAipazNdbva7kS/p6n3sGngVBvu
uYJBI3gm1llVdj+E8GwGbsREVbqdIn1k0ZExXc7h/to4+07+GMuM5Lkmhp90mh+j9NbT+PKif+9M
+CXRjXawbsnd02YvHjIYpfz5RMuDVKFgK/TauXmxUeNt5Y2+hoVensvMMgEcT8/0pjTY0pGWcmr6
yfTwTX4z/cvrtN4ZR73O9SLCKUQA4cvRFLtA1Hh+/O8dDUgWx6g/o3NmZf5p/zGw1HdIjY9k+5Pj
HYn2+yK3z2CnWJxCE9nF1meW4E2MLlvYitxxqp2pEjL9cCOMVrFzKuL5tMzlBj6eDT63CEAh4CB3
xWDCb/GwQzEx7Vq+8BfxtwcWlOMCBj45AaBhRjAOVl9pcZV8O8h2h2Vutr6qbqgOWU0JNbIq/mXO
LNU2fAig4iXioi5ydrzy4HC5hkt14J1d36KcNBVeX0Lnog8OagRVZAlEnApyQGjrh7tq4LaauXpJ
5d0GcnwyZLVNAarQ7WiGnWperRMqfsA2wVQPTn0TJBDHrV23dCBoip55U6guRBO0X0EmOdGs+LQF
Fyf3wv7fGGCAid6+4n/z2TduPen8xN8SJxXMcOvLcZaUwQk25jfyMuQu4sgnP6mHvS3DR3bu6IN/
D2NG0PGqzkivQwgaBCyHxxU3ygFhoecpB8hTa/AZy6EBLZQwiOQY+sglFPHD9Xrn91sZydN1JOYv
74RovOCvH3Olioq79iYs+By4YURXOu4YX8IQGqGxW+qBamZa9IZl5PefEwHNffhSB7vLTzaKzCm8
eHssdJpIsBeq+Yv1yDzXTxE24fJ+3JLpb2gygPthsxNojlqDE7Iby62up7fX1Vm5YTZlGLFIa30g
3YRYObPoO5pA2+3SKOdzV9jc7bVJG8S8gqr+7AvBhyDySCu36Yfu1oEFulqP9BmzqxOlv0BKnAv7
/v8yrthjHxJKK7s/zirIQHsJQJsMQyz72IOOClkJoOyUB2saayuoWlIDzkKx4n/CZ0o8Jfng8UK8
qgIG90UHSJyntZyuDCYVN/K8gyIZEevKLCDTljldVjkSxAwJwpv4Xlehn0yXulSu2xQVIWHe4cIq
1R6tUKl0u0Du9xA8jhj3kShRz64/56+dTK01XDN+bMj0FQs8GHiYLhz5ytMDpwvCl1ry9SOwvHqr
bGO/3nO0PWlXNDcBQ2Lmfdee6Iha66++AujE1M/hPlk3clTLeA9S4vtGEfWgmZdjOFBq2nvuBwf7
BTGndS+7gkOY6HuLFWP0Mmot9oepD/Ju9KsUgcQMSN09C5g7PD84zElF5mvKlzI+NMv5dcc/fYkM
wyCQF2P4q290lRF5BQNTGQysy77fAjy5/+dEPvuY+r/TRzNNc6LUBnSyEpDuMAkm97BxNgT1LO8T
2GZwxpAzTU4RKj0nXyWRi1/fev2o7QA5VPMn9Ul2gxSjHpSUOFc2mn6kELCHQJQEwsrm5fJY1xc+
cIsxSjOhdoHbYtEwHsRp95HmbiX9a5oz/RTcLJbIpr4gKn+/I3kJwQyO40SWrAoe2m9i8bt0jkVH
C3RItt3GP1onXwsJB+vUZb3lrKwAI1kVaEm8nMHHF51Fq+f+77WUOy1nr+PM5rhhWZOnKLMRZS/Q
8bVOl+PDDukDYIuvDoVCgmTYcuCk0opDaMzC8riCLvLrxEnUbbvcWLLDTne7LQtReerDtHnDimCU
+nU+gccbj4MhtBJGeBAY/l761TaujLkXdbwEzciXZHuYYA1ELDNno0Wb7O9nQDIZni2Y6xcOTWvQ
oGaG/0hw5OBOoJ4naje6107R+KFhB9BpexV+bhyfz2cSUsIANz59qwZC87HoGNzb2Axy+ojw1SGZ
iVIntZ4kKsWxWI76njm7y6nfeJ195i/CXoRQwFQrUYyw2aVDnWdrM92CGq8ebyQGgGa8AK/vlJ9g
ZiFlB58RfKE+mFXjrkHG1fFpUPH9CNzJ8BiP4SVfUFmUg7vfWFpvy23PncRsbsuMF+i2DlMBGkJA
0lUmFJR25nD87+Pnc7rpBdB9ciyFoZ5iKE8=
`protect end_protected
