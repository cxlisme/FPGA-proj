`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U3sDNM5d7jYJEIZQTnFuo64E51C+8gq0PfGADcNjuAMCEE266ZL06hQGQBM0R+DrGmrgQrq0Wrge
uPAkNN5G+g==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EY+X3Lbne3q/n8WMTQaQXRPOg34ay2XurtUPGUclFnWfBmzqnpUa8B9ymki0aidTUQYQEm2sh4CN
XOEOFCD0dbL2NgHaa05x3mCcSGq5dNxdn2t2PxrhLN9Qix/dsXnx8Dx+tcL5bK98qHkWv5TlPw9F
mQlgxUunse/mkLNp8o0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qejm1NMrPCpKtCQM6KmlkujDwbNyPltQGSiXBml/xklqOs6mwCS/d6S4AZdUpLLD3IR4u5jDDWVS
tBHBVK/11sIMg2yoMUaMj3nQivHXak00Ja3ku85yUxdiQBAhgZxAUSIYncV/h1DeR6eez1FtmUiW
k2R5zoT4kmn1ReKvyHBVXzIontFMNGOVHWDd0aaVAg2L15OVyS1Ff2rAUNHwsIDpfbkawwiEWuBY
HzkvTYgTqO3EjjRG7NHalOWEUrsKOiTJz+TKrcCeI26X/hw0q7lqif+Pw1fW7NKExvU0pb5zxe+g
dasyo7ekd1eAMBAc2D2qxnWrV/xT+mEZ2RjJIQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aEJMsL6nIvSfDKkxRVE9/86hi8XegqbQQaRNO+NCeWjYCvqPygToNaA+KX5cbTCa2ZJDNbNP0LqZ
Nf/ztarS6+Kd+yLfIhz+p4i18KkAcbPbJDi06aJfDKPZPGwgcfdAZCe9NmwjCDsNRUxF84DUxnan
NNczASRvUbnjFxV5LSeJc7fgS0ON8ZzZwIxYYN4UBE95NRZiEnndErsrJF1EiHhWW2etDqHUak7M
uJPvDNPgWyPWgFZiZqs1RYHjZsPF/LkSjAqW/s9C2dc+h1j65xJ/pXdhlNc0rO0z+LAHVHsTq/xf
4rNNAVJQPqr18LJzZvqQRta/I+LZd6EjMl3I/g==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
opiMI9un1L5qqubBM3bYmRo7L3zSLSE74WOKnJdA2zsZxyl95nt1F01km6bhA8+lOnRZr95jKUno
BVqVLm18ciDKeyCqB1ZqieL/IRXh35qDwHXUpEYaR9qYetWe96Rfmlgcs6mtV7gOqeNSetRrCEQD
RhAk8Xq9TPOwAaBY0GGCiWgPzhrabcl/GNYXx2aBQMmW0J9rLQ38Hixht17xBx15Ai50jBhhmsR0
lQD8BTlJMMD6fMBR2PAXv2wncn8avzwlLh19fU9rAxcZyfLMW/X8q1Js/JKQFdm5L0zIKmMh+rTG
91V6Q9ApkyFQcPKOXaUBzTBYujWOxjb6150fdQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V5+XqY6/KmzZKYOyYVBUe+3bN870OFCeVmp/kcSjztpDExtHlsM7vQjvaeLLq7LgsTUWchr91fDm
BcWUyxISQ6O0ukpTvBtXqh3k6jhpMYK6WWG0AxglmJ+Vrcm2v1qCLAeC6t4vatuW4PHgc4HBloHX
SA62p45b7fezLVMI/OI=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OgVTbizwEz1D5fIn9QVCVHRE9bQ/skAgyhfFYkAxhK01ppsQIEw/6DODTHQQRJeXHNFg19LWL6hn
Ruy/2+40tEWd6FxiqzXIe9DOhxqxnB9lxu1o7DXWYZWCOhfKkVKMsMlTDbTvFpYyLOkwA8aFzy19
5qWihLZMNVvFPKjEJdocORPlHzJ0Y9x0/Tlhoya7V6F7b6n9qN9zK43VZ755OaAWnh+gfIIqyyof
8C1umBq362Yld3QbRDyVlrkdxHQGPeCBFNzdyydAoDQJoNbJ9LdU5xTQJaXbQTMbdc4nayvWBA9x
Bp2aZX50ImADwqnWUo43b23foc8li+MluopNZQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 71360)
`protect data_block
XVXEjqR30uk759sv/R+ms/ekIghUDrzuYLB/Si+4+CdNiO+XRKVbw200EaYya380Nm6EDBn3oYvm
Kjr3jOYlfSrXE6sGdulUPj9LQ8TgE1Mk0Itm/s50Nwf6bLcpGewCkw9jf9w4xNYZxcoJKDfTI/2j
Tf0ILzSgLE4rvRXS0p++Ux5r7k5ZdkuouYU5H++cv9ZeZm06xTbKFfCk/5xAvAhImuNLKtffIaJS
9s2xngvHKuAWHopq1ups3z6iVQbPQDwEl8UlXZuyT2g3o8dqkpIhDg3ghqUrsThL7z1KSab4LzhS
zZBG0j1wZYgh/rzqxTsXvHRhLhw2Y5uGMKYNvhH4jJA9ozfnomvm0wTpiV9P5hzT6jJkSYlnYDIE
HJzfd/iwLNW8kYiNZ4SLJoII1i4NuY7dd6MEKpFZiubAPMBWaSndkxEFfkvStx1obBDnFC0DDjKU
YXVXhr2/8d6UCDiV2/v0KnkobEy96BcHyG6DSs8g7ONhYIolCdRfFQVt8lGBrIvSQcAG6ixlTR0A
QZLPZiPdFSLrK7+XB2bXYjebCnj8feZ7DKsTmUp7pzHvwauM4iGZxKtC933Nk9IB9I8DLnbQgO5w
qJxeqQJpm1kFll3tynqiq8vKdMCMrrHUOL0u8zDfLlxxChmA3L2GhY3idN9KdvuqkwaRYfuYXNHm
H0SCg+fJRTuvPnLOM0HlZVPGv5nKIZnHS8OUOgAg8zvfWbu3ruueFYgT8uKmmcePaKeULjwmH3Ps
tHXU4d4oGp5S4jdxNhk9Cz0RGY6KupTLlezCpGlJGSkSkR+Bhe0vIqBz9NwxKYofXIcHerA00C2g
bCjJVu1ojEsB8dzuLmutV+6h1Bqzc8E3Jgm8Y5vSMytSHEDXHYukp3oUC23xMzEyyTsXt1LvVNkL
HHShoTICuXjNTRUKMJpqaPBl+0zbBfLtfKpdSoEzQoiUonjI7knmCtBCaERNgPKRn0c4Ak5PeCIu
HUm3riqwWTfECofQo8fUFWFSMgtLTY+79//tx9z/c3tGCLObfB8LtWLHx/yswEeD7mW2cw48n/f3
9CWy54gTBFqqf6y4yAzMcI/x/c1nyWwy8nhlfGdhBSaDFZM8RMcivZakOrl7g0sZK8zlCqnZ6iwr
9gwmrjJaDlur4PPtxfAaYe84LQfvo0/qBt+GCnK5xaaDnc0RmVrJe3nmA4BOJuGQOOJkIpoq8OWH
rQSNYugrsUDfsEIHXCnd4oLnIRKlrz5HwC2HgcDxwFc/D8wLvCrtkiSpIWCllhps90hL2v7zpB0z
9KR6pwAXj7owXqw04pTWlbVofhQeEzwXDrEHc+g/LNiyNPfL7Ao/oyleTaji5ExTMYprbzDUnUfE
q7533oqZPOHMW1hKHsPcoEI/2Gjdk9284azFG3hpMPziKNyM2v4E5aGPfocE9PPeecK6dFqYxZCp
cOJjP5MeD/IsPUU18HDktSLLI2R9qHj5I5qZqM+PxQnlRKNq5CR9K1nVVzBukA458yPMza8Zo7sJ
/BnUG6A5KUs+nfiz5tAJ+GSPCG7r8dsk9qFzqc5LNF+XPYJs7Xeslxs1ND6S4ADf8hwMjHYWT6kL
KXb5Hykfm4YCWFwGKykXiUE/3e17KJyGZkYXzrXAKZ3jh8iuoAo3IU6AHgnbQa7nxYZODMMHPfkI
/65yAJFogJgQJA35eO8xYyoDkzFFPmY1q0IEka7ygREjHrrhASpi+mGWTge7k19ucZoKtfdwrZEk
NpPT3zWPH9FviGd2eR02a2PFgfpz6SJN4LNyz502x0j8dLtRFZNC0IaTsd3pi8i99HzdaOK6ywud
uwbhU++wH49avlvnVfcjURLr8P1RHDmyAk6RQKa+fVUduvDxA8tjZ9vccQwHLK6rN+ErYe0TyUQX
jC9vaKfIzGLGQJbLHWNWoaSWLYFEdPFK5x3EPm+S4pNeH04t06iZnZKlGydvpr6DAnaBp09QgUvD
VwRag5O1EyHemh3oeuvqxZBPK1qk/G0PR9jJFGiNcDnRXK0NWMrvnye4Fn/yRNwWFTaVZG0P+85D
VD7xTaSi/mymjybL7gHAq+v25IExIaTOVF7vFS17BuaN5CpAmWVrwf8vjaFfY8yaMLl0BQah3zoM
EaqWZa2g2fkA+pv6xvg6uavyRplK11sTZ9HAtTyb3EU/vGcJd9d+Hy83cJqfr4435H5+u2oGI+Y6
UpsgMOucaACROCdOAEBoVwePh+9JVloPB6k3ezs5KFQ/pKYYEfR5GfEFsNTIA1F3Fm+Y/nOXEdqD
EkUEGu1F15sjtvNLdLF/r2U7uKqu6i3wRz+hleam55EUBqohZEKmTuMbpfgy66VlJGMeH57plNTQ
7fyCOj9Ehp8j4AUwSytSgBdxMW4P1gd4mSIclJHW4IIIfJyhdex7Vy9of+ZX5PcaiFQdTf9BKbRL
rSGPAnsQSmvp2/lFdtOFMF19bi/O4Q7t1Bb+mg0hwAUfcctEg1j77Etjut9+3vVq1oYhk7wbuskf
OSUsWBVXPJHTCevy6m+pbpj37X8sbRVdaDLYJiiz2BJkPn/Nuky4KKsb/bZ55CiBkUNrG9WFkkjQ
lA9n40E5GNOXCnj9DDfp5QQ1NrnwCKsnqgUtdLxXm6GEvft4TFyL6SA5N1+VsxDsuKo167lJ4amr
EYhalHzKDE9oQrNOQNbrde2QbY38vybBE6UoyKhlYdBAc9npscURv7Mr/kmJA4d1ywDMNbdUvtiF
L4G/CbC6B2ILNijmjWqxzUBzhuJ2cPGyA9+57ljh+yLJp86eH6ps/s9sxJiq7as2SA4edGYjSNr8
M7PQPtHDSUrpy8qwq8v6fr87DOXuj7DgCuthrEPkXGaOtX4A/7JH7WUSQK0U7SuQQLrWAsw9saOj
l3O6H1kttlHZaWs+bSC8xa+MZbOnCDxXHpJ1ncakFQrqJT6TbDtC+0VIQ1dgJ0j1x9cvDVwVrNja
mStByxk/3zvrBzxAfBFizOTybT5xtuIA7gmONi87ocD9T64JOp6gbYUE2fAhqzoGTA3pzF1bTAaJ
5OykcbPCltTDkrItXU/38eWtrMjyTiIlJEOeF5icj5kaH89DL5WFTILKgtzrMqUl41VpHM5RZpVy
Q5WozIpMl1470KG8XrtgxoejTZ0zIcUfjVXvsr4hGLlVLj7vKFez3c3IOKZ72mysq8L/VPYZCM41
O/Z/GtdBOxoXwATidNotO1/0qAb+Iux9YAblHOZKMZ3LjJyU5kPQUpug/rbSDLeXJ/AtytLSeMQW
TxtRW/EZm/ITwW5kZv1Ph+RfVw4D2XKRWssNaUKk3s7Wp60Dm6OqQdBu4Op/SMpInaolpSclGUsa
ZTLyPcRlfmkbG8cbh8IcWd6B70mqDFlxQRwQP/CeREwlZkldXv3E8nT+jRmS4zNjtBoY1AwlL9DJ
7/mLktV8gxYjy19HxWt8q1MXc7ZJ7QLphg9QHA1tih20UF+t1H6l1jL8KyhMR/qhHRa2o04cieM3
dBVy0YnPFd0leprqKI+jU774HRF1dCPtS8rSFGFN9heh2cXgkiS3w1XM4oUxO/pJRARfR2nA/v2A
8fgDJtoaVEusiRfK6hRnerR5ZqFczMSFFpY+ifepve61nh8Xu6FR546zuL1o46gGQVNdCGDA+m3H
Rmdp1eZji9rLiYKIaQOTBc3hQbhZaxJkmmIxKAimjToY8Byjv9js8PjzFr9B22b0V0YFbu4sO+Nz
iX02+JOJF4BSGRyAPXr+l1Uz+6zdKvw2pem3KYHn2utSJ4BMWoRERK2G69pOVHmfdDkvbEkcfMaM
udnBAiRN0Tj1Ckg2wOjk3lXwhJGkngLAvD9obO+CF485tGKh/WB8yO37Zs9G9orjqEcoFJho20z3
s/TgPDjlbuUZSgzxD6uOgfwE880zvbvDukKyW41sjetWOoRiT1NYu4FY5+HIRs5D/mi9/1V3V/H7
Tnhx+aD5P6yKcNwGgOOdwa1h+kyNi2gkIM9r0B6sYK+mm/kj9y97FXZQ3gBfgwUO0mb1rYyLAovB
gv6rrZTBVXo/JlFNq/e9BGJF3uzwCsaxFDy4TXx0k3DiM5TMlJmlj+kzslL/z+qBq93os9LZ50Ri
8RBirjdNymA1X+SQ/6geyUa2X6J/kGClruyl3F49ZKJJKO6Kf2GHLFbtj0n0rpiqukmSAkF7whHE
LioniKj1GRp+RoGsvKKEbv5dFFfMPO40Tl81ivz0DYHup+WeoM7WF+XVTkW6k5jFRvZWU5O+CYEy
cMm/3Ee+X2ZaD2wRHoZAeBOOZr7USOdwdWrFoYiFkAlfYsqid+4lce2XsRwm47851FxridbvTnew
mKfSRc3DcR8BPbCFaqAR8ZeKjKsNhR9aDNu9m3t1nwqMrjuAqdaF6j9ajrV9UfCmwS2NxXS8vDGU
Qy6wLIr+iTjMGC+XDil0z7emwMDdT30B0sIYpsmrcpE0hlwMc7hvANzlNxdUez9TmxWGJYRTx0NY
NrzLeIEczLcrZKEqEJGXhOXkPrAdR7g6/KpRC25OnE6ALIcLCH9wNV0cARV+Nl0XLVV4FTpk++Co
ZbxmJeRp6fLfB+boPWztEq204us0KzqXccBpRDVJqWgEqvzhgBZvXgiy13Tr0A4/jOCBK4Ac31nO
insfu15Cc7LqHCbingGp6xgWxa3DRyVtnP9fAW0xQVLstoqK1P7VlYbajmNiz6x6/FASXFA7pcIK
1U4usu8Q/uVFvF5IRLDtdJmYWKuBw629fybUazAHdrY6YhNAkVh0cbZn54gmF4ixqd2whv6pLETU
MUbOAHWQEYfCx416m3yfTrjOX+R/RdzzlUA5LjZWJrR3mt15gZBL79KPa/2w2OSKWcQeWGoCnt7X
zYGGevyfSfpvxrffezGIMQPswR14vVjq/9zpnzPNHpxWftQhgUM5dYcCZbx3YuOxdI+OXD3IVIXT
habAQvN2gGLsSx4/aqm/SARubFcxv7YGLtpaxVnmtWS7AKsxoJiurQlnHO5DhfcDNGXMY4WnIUPr
Y8wREkSB0nHBNJbALyDdp0JDxa5jAVB1exbWyH/BHr5tVr17i/de+MVL+is+kpDnWwL/09AEZpG3
8tXGFwgZVeueqTcAtogJmZZ7ujhi7+f2Axx9VH9FCT5vD1e3PSrGKTSq1/MQYqz+RSQFY26a9Q0t
S2kWiBs6ZQDb+URDfEWwMVbeoVxBZ7WzQJKKrmqG4TlBS5fZMBUPzBC7cqX1l4gLlEo90nwT8GSn
DDQL8W6r8e0f1Tw9/OrKSWWgwGmFyBdYdKhOHLddMqi3gGwDz7YQIfEk4OhyzGr4en/046SVcXlh
SpESrXiM2RHXYxjSqspr/PqqMfhJqAxLHCPEzGhVvM7m9yy9a29ZJWsn8K5HUwmFgP/AOMLbqsTE
m713YMTyLNgQ+rHRjH/Rx7L18afSIjjZ/4nyhkCAn+IB8N7G2m2bsW6AfrpcbrasJbFRdkyfAbkA
5YIB4HJLLh5TSAYuOGy7RaeyltSMoOgnMUbXfAWKX1/SrR4RQN1xjMSnJ8H/I6GdlUoM+faLpMY3
jNXHANrV92JmpZb1fE+KSJhsykeE8ULk+E028PlFr473wLdgLTzBpiwK/N+a3NDNZ4piS7f0kVVZ
Yjx7Wd3nHXWbPlTv+pDkgSEeGMDK5LxYlnvsIy9iSeROIrF6xIt2TEvF9XVi1/ZSncilpuOC7ah3
56aJA8tr4YuHjkccvOQd4wTISc8/vpExtfdOdJaaf7oCfm9nreyAU40WptQKY9UcTDjIzA/VlOYu
c8J+iEGR8VJ0MUiQTKpZX4FDFuCn8WiKrUFaLmsedO3w2OC8PCUJ+SRUFXlchTZPOtXtq7CXeIde
0B/ym2s7SqqWwr8ObEtOhCabSr/koKQrjZJ7H0nmLvK4nsBgUoXlX2qj/1f0B3R/kWs8QxRF3wOz
t13l0sTqvrTgaC1nLndf+YD/POWUIt53svCeA/9uZOU1zWeYS2oS9dOSlhgDDeEBajO/0fl0YuMw
N05S7wxYhGT/CnPzCnd0pzwz44HTQqwqUhJv610nyloFMldhsIy8WGVw1dgwVj7TvQniXOdYMJUc
oDj7WyNwE4LrUxnwqgbQOdjb37ryRhOviCW0AeKuP2wKsaU5fE44geJ0nElTuPyGjEOfVmEgvx6V
awEm84k0XPdbQIQmcToeStR7kY9hzm9mb8zHNP+8IY8vlaJw7jYpNPYB4HIdVK1I/y6qSiqqWMz4
XiCk2CQ7nTlCbv+7tm+i8G7T1vNAOu12Sgms0SG80tVeInmR2I4PgHKyUeErVgffnnokIRzdVt/u
sX47fhEQkDHU/JSCJL8rJTiFlkg1VQ7zheYWmMulCVvH8UdlKyWeuWy1sy5iRu6bIvYuydM7PAlP
fsQENpnY76MzDiiSXOy0+gR9TI38fCsjrRubyDxTQEQf7KIzRFCQ/YV2b1UFjrz8QhFgVn3fb1a0
QP2Ei77cUMp5EpTT58icM3wpoU5xbEpcLGMIdohLtDJhazBhpoQjgSMSiLKd2ayoZsVbV+Dxh889
RaHuPbAFwosMY3uR1pA0A/dB1qPEv/gHzpz+4LdKMi7Nt3gmH/m86Jz7k5nB0WKUkw5Yubhj2aga
F0gLg9nxbIp6DTrhYa9gJA/ExBUC645hgGlCH06PkxFWq7E3mkuRn/3E4KyL0vD73h7B72QC8bjl
5XY7jdcckIY5yunLJHwbx9JXJxVerrvdSnndGyA7aekTawR1Ei04y0lJHtyCosEwjtgMc7s0TFj3
37RWE7Rvk9SwcRKSVAVkxQDj7nTKoQtD6eoLlkbu1vLUKAZbVMtT4pt5qMps18uBs9xMjW0Eepwr
hXYyDPhda/wO+cS0C5agkfQRkQ6R3cK6r7c56Ot6+0tRvZQOGky7+RRFY5pF6Ayk6hRmawziHwRU
Co1FrhnQRSuSLRu07RhedIkCPOtB4TzOGRAqVuJgrUEW420cGYrHMetaINNzdZDAlYCVT8d4BK0B
J6Mzu8QTSgh7F/ng07vj5/8ArEqy3p0YenhY/7M/Z+BOSsQoAa+9O48eLwVEho5icIX+I5OJsaeS
qI3Y7WImct971b1clgM8G8susacDjzAGXAVJTB6+6KI09lgLiRBfaeG20owyD/7ck92TawBpNWC+
7wqn/iGZwZ2WcUQ4v+/DU/CCDFb2DV733JAvfa8gysmBDR/Bt0wILQnK3R3s0VKCRtIkvn3FNHiy
ntCdkkRd1fZAcb58huMvZ80qL3YOD069fAxb0PZkRG3umeqHaOUg0QihhwTHHpcql0YHwKVp67cs
ZS1uOMSpxHWuxLaOROvLCaVXZ7ATrRXJ7tuOS5sOwxDTBICZ7dKgc9wh+pWuHiJyE6eXOXlnLPQF
lG2EQ/sOH1L8YlWkBOUgIfvWCHVn7FJTF/rpe5jzviql/CGybZZTACnrLMBy5czc/5W2CkmQ/l8j
eJ50wc5LTU7NagweE/41YkaQQqppq0B8laxWuo4sbYTRwjDzWggUDoVs++2q9LCpMq6/v1v/Wd5Q
PlFdOzO49sI180CAWVUFWzwRnq0FhgbxjQujsKoLEQbHQHjXBzgkthHKgWDXSayjNZDeVAfNCi/y
F7OPXAtFskPTccxF9knWkLzrRQnbYbUV80YxfiWX/KAwJW5wiS09YPaDgur9Bvt3A1Z6BfGfJFWN
yjX1IoByQ/FToZwG/igObY9SLohl4FdhJHX4EGAXOi2H6fEOPs700JacZfjCTlUy9hMZhZx7xQvX
L8e0OTPMVps5NNy0XTS+N4Ar+EQJTOkasQMSexnlmwTPshAAXcuxXmg4NjZ/7he24C+rthRnE1X1
msq6bGIt7C3BsWEP0lD4gRfyV+kE5QQiQNjHSdMOv2KJVvAhibgmLUvoZgPC4kdNh2HYC/JqyZLY
W+FwYzEINA0i0Gjx/or+KRI1+ceI+CCjxVOaVJ4e0KaT93U87zqnmUB61WxSlAn0cXY2u7u7X8Di
olmMq3qkAJidnkzVHbkNVmGRjUdfJa37R+SCs+uUGb3HocNhv0gmBV4YDm31/CJDPY01tr5FGG1J
sKR5CYzwDpFExbQDpRd2PBOYkqAYF9vV6Ft1LXZjYzJeBYNC59YRrDhgfKq+MGAniGRI2I+i2pr1
94UFBz+0LVhttPOYs0U3Qqt01ePboZKQOWrsIfPp400EfF5nButcN4lGmf48YZUkXXMzOHGZ13Qi
0o9yOo2b6ZOnoQDkstCV7hSZB3r+9ByGFIEs6c2c9+UggRb2bhAP5hAwPduojMuWegGW9oqBP63g
c3tVEFlm9K3PG2wf6vTCjsw2kmNair+5OWRdKj1WBtewP6vwHwOfLqiizIrd8Q2JZ0KGLbcrt8GY
C8J+I2SPupic1ZV2xNayfexb5+kTN7YYwMY4vwZcFfqUK3EBUN2oPf8F+lJPc07nraayu77Y+dzJ
inrBQmGyArvcow8mWrjXMt0mqBMVlMuMdcyvARYXxfnBOm6pg2EmSRXjx5m9eftWdtpEoNE1ou9Q
ibxGLGTQbBNqGM5wR6nnmYCESgzAD1qOE0fSQoMQZ43xHS/J4gLwgN5ifw30aqNRbd7DMqEergQd
GgnXV3IwQpyS0rIlEFAnwecSPX8a+L0AMF98b5JGRiqe8RBvFr4cF1ZCK0Epz04YEkQh759T6sPs
vbZLr/q1CjxjxRUgom18JkT3y3Lm0WXR8jKn4mDViGEt9FElEJCzSi2fg7yCk2agEPe34nWQ2+bQ
1apF+2vM//q7yksD3PBisjHfMaPM8i2F3+M6Uk522nxQ1qOGGZ9yRjILtmh4Ok98+opCFed1WBO6
1B/gW9ThEZdL1IjIBJAskrehYl93MO67+Xetoq7z+W7nBLFrWctF8hI74uzf64cPc1pnNFNlIS4p
oI6s+GZ0XZ4tEDpCGQ3+ThBHYvA9zlxqfF/RWl72Mf+7EJYaBZWd2WH+BqnpyFQKRKZ9ttACW0/a
J0nHaJF6SCBPF4v1yDKyu8c0TsCCJ+B2Lb42ySHEaRKtzF6ZmZx7dngcdGPaWR+lflxJzjJ6oXgl
ZY3num3tIi/v0OWVSPkCHx/nkEXvVp0NoUjjL6czaZWVlFwaIlTEm4ys4oCS4HOn0s38G9U9wpuC
WQ7265Nww90YsisK6HsuoHeMXd1+eZk0iEw+35cac5xT3LYo2pck/rt4XhnjW9VxE6slt++O+QBN
Dwy7e9xT7P9f4hRLZyNWosOsokCHYl2KrcRKeQNuP0UGZVdKbd2cyDmSFqxwIXXzSEvVbAePlUGW
Lrvb9OlMODr0pxieK9ebNJNIt/F7xUUw5Ef3roHu+ObQfE2sczDjsOgK3fMskCRG1FCyTufrVkbR
pN3Pq1+iOMOWLADOsGsF+a90IBFf4pM0qyL3/z3Z4XiDu/43hJdKIRSgkF7TPh0sKAqqR2QGsMbg
aI/As60sXTh+RSCm36eMv2UfrF0I+Ivhjfv6QLf+7vuNpddFFKeO54bd84bTo9gtStvo8Rw3Z1la
CD1tLgaPdMeg5PmWP9vR5H5X1V/tfOgMFf3Xrh7ec5sDlXPSG6FQtDlbW97MNxzHaADVtlwTGdKm
cI17UlMTvgp/SIjIn2R9aZYwTNlRhJvGFS77hdFQBHc7l/EnExQRAoyiJX6OEY4UCA/l6doYD/yS
JNN8tfUQLIZbms5tn9FGsfxrF7C8HuFiD2Y81N1svO8X2y5mkML+YnCAcK5kCBkqMi286VaTXTuW
iJ6Fq1H2d+0WLDgHjsJFSz4SGylLP10MIWhf5K/uB9p+W2oie+zyZzAzM2tIud+17OkqEafP2032
2M5yMnVOwYmDqYmtNmKzvbIRSeJvt1XMOBnMJoXgaZYWR/cyJ2WcXu/ORVq2Ur1ReAWSSWV1Ir2j
6qTZDXQI64gun+9elotX/HmqPKzQcxyoSRo4vshUkMYANgZYXLT1CRhZct0iMhsjQU/hmphDK0Mp
Iw7cCYRvvGK9CJAOKldkUqoJAlHMqwLrou9y451fPUioq5+1n1ScWxzYoqO9mnglBc65IyeYjksv
fe/m/ewmfGO24hRoTSM9Pr0pK4dxmWO68ROMyWwXzTXGOPDwKk/UAJzNIP+M/IsEe+Ju+gaiFB7m
U7M1yI4SHsk7t39FV4OExN2DwlE66wYT0iYBzDVPmgDx+MswdivIRleDoaSvTQeH9cS4d6bK5vtU
TJ5zZBgeb6qs9Y8ZrNDAoLVcQYyKfvd5UhlTvPI7iFbGhUWupZJOizWR3mqKQQph8gFadQ8QTjjP
77z7PnKbncSK31pfw7VOcAkjwZBLb3XqWq6HK06Ff6C8L9Zm7mZy9BkfN6ybdKRiBiFVHaJK7EdR
A9nBGVcougnb2Rzf+jC9RFdkjHBMXv4HOiGmDLK3MEWTLNeWxdWQctlL2sm3ZA5xA5VoJW98M3JZ
RF9ejdG9SWO6zT449q9DEmU5AhUtWyyD1mib11LJxvx5fgGahtIUxJ/PWdUh+KLOeSsBTpTYuVdR
IeN8EzWwuCdYnIuy1YUn/Z5mvu9df1scccfOIFbzHCgGAA28+W0/jdkmHJBBS+plnkFFLk1Ac3/d
1fekDg0iWu5cg3UhABgSwoL7ZpM4BzlBVJmiYj7KRWg7i1obD1FmUradIdeoPlswD0gBmMrWeUbL
o2rHoBHKY9NapnFX8+YAIMe4P+6TKpHskHB9xlDvwBHVFdostCuPYBXrSyh1WB2ToJYZWCT2FnB3
FzNCg7Z94LEwZBNh+/Ztm2g7nYwEnwHugu9l+oGSvELTjAzZ0WYNDBohL8seFkS1+x611lB4RPjW
vUpTPG/DDiw3yVCFAwuS+3nrFVRYXbUqhM1xiQ0TliktdhRDnTUamLIOmdZlOjDUIcsh+1KDpAo1
lfhnBiIt3SEd0rVykgXnDiYXxpeeg5DlvJmTxixfRwIKs1fkUpo7WxPznxo+JOo1Dcyz1d8iURvx
RPkhJRqW9MUYJgffxGi1m++q3U2h1HvMC6c4Noonrnl5Ml+QaTDf1VAkOyA+dicEUKXN7EcDmnbm
hV83Lee67bb+IveUsxQvO+D73DoFwmgWK8aMR/pzk0osc1pSK1+pWwBVJ4qu37epf6aOwOPOTXQr
nUnJD4VmstmbmXxrhbNIT3l9chv4UI8xmlkGzJnLfYp7eT53YzcGuhTnLUFSuJcSzeEb1fJz/eST
Xqk7fWWb6X6Uyi5Vb0DTyit9DTDyaw0A8zSfKgnAYHCHg9ObJdO1Xaacx4o7hl56wMTZttM3A2M1
FHTPXL4Ny4Hk33R3FC9dKeL+nAffz96wDF9yDExYN7BvCvO5wzLzltMi4+2aDsgC1tg/19dWkPXw
6eYMF0MQTH6WfB54uQKc3Qf2idQ6Ksj1CCRECgDE+pqHqDNOkIxoTMITvdjl0Cw47pSbiAmYga4C
WkARM5lbr8iUms2HrRb7b5qipyKsPSxm9Nvwz+gq0lmm8RpNHRowHGRZ2YKF9+je+zDY6GD9TbUu
e7uIIwnF+waDTtpPmTSczqpa5IrgDgPeajRHzmzFYt6ZTVOxX2BlieG7sKX7Nolw5ta874he4jY9
YUwps1GVT6Md7mxgtLbmmOOA8+lmQTE4wfcu1yfZj2HeP8AKRF2zLMrO32cdd4jdzmKgNFHJ5eXm
JQvLu8+6L7m6gODMUXgE9eZLyospy3TbCfIlwRVXPnRg9UY1h/hMpZ0sNmNzbLJacHxtPBopYi2J
XbXnOwvVgWh/qZrtbuBIkQVs3ibOThTHA5VvVk4ThbmhCVCceK3w4exXDKeRRFQjpE3HfwhXCw8m
yNI6hr6jgUlXoR2IaAgEti+ouyrZkiTvUIpdAReVCuEvdCkqiMQ7IDz+BHTZTXF+EX+TwuS3mQ6J
E5LziEjCDUWINw5geOQNEJfVOUwx6Aou9/zfiFtAVXSPA3zZG6FGs6dltGzq2i8BOSsZNvYelE37
7BLbaGdD8m4Du2SCFRr2qM1rOXHad1Ql1MazUn+cVhPnTN80PVNeAwBSRavV+u9RSmOIMsm4kPWO
/5kaXbUUNwFbk9T21V3CMAak5mhlNQf4FH7ZqCtvVob+/t82ZmvFAO4ME7weTI59G2KPOB/lIw3c
Z84TQMi4yn7MD/9GA3537oWxDcXvdqg/3CyIeXdQrFLwJNStScofdYUe+1D/y4/+pdGk4dfHHkIw
tPMYHUYPfFejdNZIcE5gkBfoyGHNBYs0hJQGMKFo8Xv3yEgX1p+Dqkw01hgtRulq41x04dXR82yJ
3k6LB7TNM7Ubddx1+o9Wfad8oxHHvkx5+Y70d2nNBWI2aFcV6tq9m659jY6UXUMxXQ0BK/JhRd9b
mILrOo5BPtHUG1hGG/fS0/2SvsYeOWDv6PV3LchfbuZlK1z+sjztPa7HeH/NRGAv6C4QoxQ1mpw5
uUygcfqfb2qvELJfqcxRBLEtLDuRjFvq5kcEn3rBKf460yT0Cjas4KnySTISSvFsDhvGGyciw6iu
Q6VS/B2r/ym6cskPpgLgR30PL5k7Ibfmwj8OjJyJXao+ervY8RCBwcdB7eGGCtsbznpeNhTEQ350
06KGnhlJPP5XgbLMXrcv3p5iZhOS6sxum1Naxz4xUQa7Tor6gLC5P3zZsViXBebfwVj12TksEXRc
GR9exVcq7iHJmyPzf31Ba87ac/woq4kwverrSzYlhfanSzHN4Lya+UiCDaWWw9UvMJ8bxSOZEc8O
d8wW9rIJPck15UlYnR745BNTkxvFlhTxyMl3oh0VWTJRXAsKRzQTDkjSFEC8EgabS2Cu4IM5fXY7
HmLCTtSoLjaOBk48wLBMKYNuASGvszlPVX3D6EFADlNJeRSwz1pk7Lad2zdEH1/c+AS4DJegyIIg
LXHy3TXqyNsYVqtUgFdULNYb5xJLISb+Ka8uD+4Y9CF/kDm7ui+4UiTYkYIt3WgF2DMkJeDcXK5X
d6Ks9ZofXYdR5qOGzO1GTD8nhtVHPz6mFOKFhd1qUOilF6oR8LL1dLm1+hquI6q8zvrFfYCHKAuD
Aulimu6zQJktwJS4QgbwD406n5rY/w0PWl9P/uXl/83FbS2UQ8VRKbrRB9U7ZB87OEZId0MLHywT
my2c5ydkwsTMjdpUb/F5j2fqk1hmXHS/EBOCiP1a2+H3lHoKKSl8H38ap1aRsiEBK1vk+pHmO/yE
/mXWFkGA1enOgeCOSXO3bbpMLfwKuPw62qlUDmFKSpYNfINrgLUfG6ghadbOpUd2A9TZI3p03DDy
/AYOf8qRd+NrK5yGSqbYHwQPmzvEgrXCZP/bHDV8QjWAsli3w+zxKW1Wb+hnisbkwxepcRgH0g4c
nEdTHL/iuebh8G3Da1hH/X0LrVbnkLw5aW7SWa5zCNCWxtGHN+YwQOfe9qBg3pgy8VCObzzDPNMV
BQwd65mBGn9nXhbwdxGIDNF9vfJfQJ3uObhXE/dqttkhGjVoEFfQ8o+vvpbDlnteDZyG1+M/uEQb
EED27GdId5JmdICwX8tCqGoXb6sQv00XFMBE/MFMMJmdlvltuZrFWPv/VFm2IXD8rQaUvy1cIpfT
J1/M+KdKdqYuok3TpEpeb8BvUI/pn2t++m/L9u1FyLfYZYsmNGpnk1dJDjpfRmD8lENGpdo56NtC
gEEUg2z20qF3E0sZCnpum+gQJ6XgGK/2ExeczNpam8+nfzfu/0Eyr7m/YFYknSMoENGYacFxdLH+
DW3kCJXSXs/JV/9Oh5nTgXMKF3Z/WnY5fcL1QYAKeYrbJ0IWiIOCNW2uX83vNUpVGD/cVrzzEu8V
z1tw5w2Q1uQJGgJMqKhfKj2cuO7T2cdC+VVO/AjqzSPaRnsU1tlaAzrbrgw+a7hlEh2epBFUnZ6l
tQG207X8auWXAKMzJlXzCwZvq+I+Du5+PYsS6hFn7v5rE43v+EZHCqf7cPHh7VOTcXTEBN9/Aqcc
2k6ATz20g0YU25VwFtGztSa2pqLeByYiXU8MF5R4rsN6sg4ss2/s683AmOL6XGP8AQw3QdrbDnrT
iXCHwf+CHz0FFzyzrZ2DNCevWGbs1XWMH5O7Vdf1USxOa5rJEEahBpB3e3H9na68riQq3Ut13BKI
FEsQTSdrxWPv1ZtC3AOLCPwREGl72Nyrn118YwAIcfIci4VwLwyHZ4gDLKrNCnqJWg9Qpz7/RmxT
Mf8qjVQzukqmsh55wevj9XDTkTEO0T6Z0QFNSyLuwCuKn6tolMpWdIZRm+7G5Baxa7JPXmTM7jbb
SYRGjpqPeuw/PNyl36vC5CDWnoW5wB+2MteFDYgNF+WAk90e7A8ABm9jjtWwzJohEejxZo8B/Yub
CtDpqqOjoL6maGce1MXvm+VGZfsO/aeIH1lIpI4qiStfPTG3wgNGCJg/vOxl1kw+DcCOnpNYP6KK
ySPDnDEzyz5Y9C4RuNSMh/UK5tHNAKnIEnx/dR63nyjzwe091D74D8xj1+IZC4ZV9HurDaq8uMpj
Sb63edvHBOgfq1e3eSKX/R3yYIfAAk2BSz2aw4ujM6flsxNWk4WrwPMZd1OwZgfa7dIB7QVM+zgc
LXrdYioyFB63/Ehd2y8CxajbQzOHVeoPbXUHmLNTz8pZ+VGoG/pwBR9q1DEZ377DaL+q14iImBvB
3BH8mCeGTt06PV3jMb9UKxZ9jeX0njTCdEQoQSP7Q6Tv7RgkJ9clSLrBXCvWCIkxUlVBVKUB4t9N
h5bZzQ6BZ+mT96RNkdaFXWpXPNWRY8oi1L1yB7ePM3N+olZAymXLqA7OoCLivZrUmidEuNTU+OfZ
klfZ7FQ8Z98uNUFbvsopqoj/dkKA0YEPDKeuoKQcFgcZHWVBtJm05p3vgIGZTYF9Sn/lr5Yb1dgY
AY9Q/VP6qwxDNTEokbxPRZmzmyUlIpuRuv3WaslnSqwjU6n/rT0OyYuOzgbH50/wmlSfcLPSk1v6
CIRX3EC3K/ENi9xahpBbE8Xn5oDdYqNrkoixhm5+ErHmVO1RhTlZXKVDfQIXR/P95H9CTy3lx71E
1aMcK4KTTxWpyO4tyrFjtMB//bcu+Q4Lg0KaSpJhpNWlqGAJv6+VOYnxdieEv3V8WRBBEG3a7bWk
RmH4rkRDwm0iLq7dPNvdCF3gbEfZ90KsVQDE/hiZR7TSSrukeeAsuecD8w9jd/OD7krpOwC+bzti
mViNaFANrWOgzsn3hVPgIRmCD7OAk2RQSFCz8fIqwgmgvYlCWgGKNY/v570p6XPHd8hossxILw9C
E+JZ0rDmoCJCZQ1If2J8aueUNuze1zdKvT1CgxjlMm+zFLoM8PDfJy1rqngyPGaNM97YHPFpX5WQ
2I+YtUXrtHio3J/TCY5SyWELix+knYEsfbhzOBv9eHO3DDqcuDGjuplpcxVji8jaCYy0Tt9M40lJ
vK7ieyf4TZqbA/xQMq3td/W3umdqdfIbWmCfNYjsUq3u2adBbhDGIQOBM9L4SNN71/dv9E7iJ+/j
941fiX0K5v16bpcNQFJnKuy64raijULQC8UfDJ+rBd//RBX6mCLM+25vYFuGcOfON+Rmdc4X1xLs
/qW0nV9/3dfmn1Z4R4UQVIjSJrXZRDhS1y0ZQwErNnJ+jPqaczvaqPzWLFdxz2KlXDhn31K8HD5O
VqChh+5Dvem82EOhX9kSmzRuee6AF/CnBRidqdRS2dlT1jta32POSp62nhg39QfsV5UDEgB5zKLt
fHqWazHfHCqEBnDAGlmqyG7IIBwOgRQ/46cMAIT8TYtwP7CpHhzN+ybExcej+9J3UEpLksl/bSUy
skQFMudbxY5Dmry51qilrKYYG44SLV4h2SIjo1HfWTAKhr94Bczt/TMljASZomAfx19mUSXXNmGt
lL+m6RnD6rTWQSXehnIzeC+Cy/4f+7J9Vs1N9G8Aa0U7HKbPegQRK3lt3d1MiAJDjkpPPqz40zBD
Uyk2ukX4puKIELKtkPH5ar7JGTyE6mXlqEEg9g7qv+7oTTNayg8FGwm1oOehQVX65Ic38Fw7MnX8
V8/FsNuM3VCnRYClS1WPeGleMHScnYlZnRpY91eqMREn8wFW08UBLUyitjsC3raFX20tcnF2FDiz
vZ7OfJdnHdsYD58lePPzaFYOtFpxdzX504cV8LmRoCIj/G3izlxZpqnZKlqszShtr81Yfa29PuGH
qxCh40+Uu13XR6BH0nBHvAGqEJs/TnMpBgU5ExLtVdeY9/GEBX4ue9x7zMZ80bpdwAIwZexANfR4
kJSgJp9bnrbQlsbWUPHGso0GJkLoZcjOC5t3P9YMTKWlcX+HUGX7ftOfRfhQ5fXNvrFiop2Kqa6j
H17FH+db5BFxv6MNJUrkUnZAuk0bBecT8OST/xi5D9oKjLQsyQ1PbR3e82uoNEn2BSN9dl7MfKd8
oI15zcGQ0sIzP/PZ1VlNG1t1rZgOAF9CTv6CU1sIvjQ6Z6TXOrxi9FKCDrKFReV3dSt9pXlO2+f/
n5OevIY9SHHp/7LkeLQ10JUM4LoQxjSpcFP4FpuzAAtbzVectsFXSGTnjbglv+14Wn8zHkNE4/Oh
SCUSQXWoBAdUHHeinOWM35OYNSRU8BZ5ghxoLRD5H3xFFbG8N3QVUxKswtX2OGp2WucHteDHmP/k
EgGYn2lD6DTNv/fVSlx/OemvzEZGowBDJ1yuK88I+S7VMlmRhB5d4XEZU+exaO2Y6b3EkmSGFjYf
AIRnF0Ty2wH/sIvfli0uWlA3pr1bZhTk6GL+ZHbBA+p6cIc+HTXRetelgb7yOHvqbOqaxKtniYXj
GchunN7Ovuoj2WCFkJyEWZ6QNKX1ZN4f1T//A4ac1q58VJryDplQcnckKHJ49JOCPlv1DGJDw1Iu
O1p9lIlHis5PjZg6akmQqhLyS7Wop9j5ylbw3lGIwbzybmtiYtUaogrjx8vAeiCBnBpCiKOt0IBL
skf5EcGHqB80KYxMLSqHIJKI3/s617Z10ay3O1wnUrp0hni2L7n+4PIOmQT2ui/axkVErmThMiMe
1QOxwTSFOcdaOdZLK8ahziY1F3KkiHaa3djliQmYgJCGqGTFJ+wfzXHPPKDDwl7dUT6lUJEIVdOp
KYpEih5WYaln+rtI/8gFS4XrfPmht0KOWWPy/uX9LH+dS/47U9smQCBK5ayTplYRe8UYlbFs/2HS
WyDEWEq4DUWGJC5EnLVWM2GjEMlDjc/yg1njDRTZV1dPoDvgp7dZFN4bf6adu7RyG381uIPsLeZr
Unj7WSTethtMZZgTVqHAjZM6XWGMuGLhbdc5QzaGUBFAwnsHd1R9PotGej2bIbsc0s7JMPf+oQrh
rNOpA6W14K1FY5Gd+/VXJXZy/duwifI5VFUaO3MKLd4J3EmreT7X1gbClAAclbIEy1RZzg+zzZfe
DL8NecFTzg/m48d+TMNtbINm64TQRU8gJjSwPOIjdAh8HeQB+g2jV0n8/aBJESSU9t6/upQpo4Cn
3Ht7dP1QZ32Ee+afHFOz4A3MgC+Wzex1NfkOiTC3Mv6vbcYHcSBZEKm/qd65sReLHpifSvaJkJdy
GdhQUeBh5l4METFMXvo/mO50fuOBG8hNHlyNkhECQcE/FI+n0FYDfiGGtkbKgiXRhID9TJg+QPbH
aVjnwSqpxZbkUoU9amoP0wYlFAt31wfk52m9wNkGbjKYPVso1gZYY9bHlOjg19M2flfJrRT+X3lI
NxuCSagv76kFsFEMKvz8QceMTY7GwKMV4/J22SY6CBSsN/bmKsY9W3oSCFKvgXpLotCD1Bhc58rc
lIGvgprHIbMQ6Jlzp097yttr1YWWz9EzpbciaYFc4Ytod+CvIMItNntBCdV00jWH4MgeaZlS7hmx
UbMbr87NWH8svP3/D3W7MUo+2ABLh4NklaLO929EPrM6EKLeGgvSb01dRjvoEuXuJKJy/QWAcFSt
KO4RMTgG6WN6Gxg+NXhEs8CLwnQbCO96FM/x24cNrIba5fibuCau/qTcVxmd/Rmb+ZWNAvK/9HlO
qZWsDVebuL6PCBb2qMEnbtW0AyMkB43zMwAEaVXFkYE/8I1kZWhwi96x5tucz5ccAKW1tM0hfCDm
L9y3N9+ZnfpBIdl4bC3fD6DJWYuCXrEz2JyQFWvWUucoKwzbGDyyE9GpbPyg2+SenH6ahLMOeFc0
qdF/dVWvtu/yZJS40AXTZ08ExV/LwgkRhMx2Y48SB6I2D28ZwRuZ2n8RDB4lo5LOI4TG1JsoTHDd
9+njB7WdKLLBR59qwBV9BPMgcUApjVickfZEIl5vlibjmUQQ5ocFzAiTWckAeTWvegR+4cgYqhXC
1vqdFXivH8zuRmF/xQxlm6K+qalOlsdDAjSDwl5QIN0OXDkuiZhY2bPegLzqn+14A5op4GJaqXsD
8ukyAedtQd3lLWtyQsHVcDxT2O6LPAT4iXXrvALe9eEj4NnqkKFHqcBH7I2mvrAhVmzKER834k4V
W7pLmzQQQk1MOp/9YlPaSUJpHbTqLkT2SzQoNxeXH+J5q9QXrKdXDRnWISgg6MfTPzqnTQkIGAeQ
/tdP2Qdm9J7rBAbkhCsu5s54b0IIXWYV3NCH3yasMhBfis4wneGuKagUZCSmk3gMBP7B2+qg7+ZT
zkoCQP44nxiLT+CyAdE1K2gOZVfzsy8TsqCtKcrcp6yTn6pR9Pk5BOs/T5n7ZcXk8iggI5qO8rll
87pRmOHEeuofpnXlIlafVXvIkqpRWikaZU77Tlw8fWaxwqjBe4EOjyuFV+mv8axp3zD673aybuU1
EGiYiwNHsyHxaLUd8g3NCGngFPO0EnvqkAyJT0dbPrW/TQqBJYehWtbGlh4CH2Sf9qH6Mn2WvuqA
tRmp7Cp3oewRrWV52d9tZcEkk54sLdLViLa1+4YE+fMW37Z/gbZwGLTa4JAx2ibRYvHbAbvt8eLr
e3gEBxuqoe0zL0KFDA+D4Hag0oyKUzwRBDhbZPTarCl5t3oXd2qP7d/gl7+PtHyzTaN/qJ2SfNGv
5sjigViW0or2wLU9AvArxcdsa/0vLIiP+Au/JClIMbDEczCRZvI+ym8AsV8FigByL3yC5EvKfEcW
UTNlm5HCR9sLCB7kOGU8JbW1cRI3sa0zA6yWiKj/Y4zxInxXQ0FhAMvv0ZrqO35MNaSu6xeE7/bv
8BQ9JkwFNOwq4JrmXeiFANQ/Y0RLSGBFSX99dM2m92JRmmPinikkuQaqZoZIpJBtOJWdpJvrVELW
R/4OuB9G0jPhrRTdz5MhaqhqKMSwrI8GR4kMUKg2P/L0p43SdSn9619txfay6WXCrdBnsXnBsmE0
0sdqKGBrdbsOim+ApSuGfBpzU7gYH9XQgmJdRLVsnCCe1pgtyEv2TcFNwYIPpjupExNSq95zKzEC
3g+S+x5myTUTdUGZjTynQ7KojYJ7VwPhiYKuesnIi6avt1EfUxTAOyO/r1+mXrwTXVTzWG5I7YMx
nZ4w7z20o0Xn6kLD0qtuiGjIHZg8kSIHhjy9+MCkk2O/6k4+QR7fFBKE48d7KXkGGclBNuRRAbRT
Mh+iYZFz8f2it6aV11iYrWrSw0ysbhUSHj6m+gXLob+UdZP+xgnsMIslgwWgnnTgoe7Cv6ETJC06
l6TYvhg/hQ78UaZ6ih21bgWLfzQWJSeqJa2Qn9duCA4iqemOm6IaP3ZY0HUn8+bQgoPF5r1s1GbC
SztL5AiJS0eT48sh0XqObkWIDZgVt1OOhBDyGcezYEr4CqIQrsK00d5GyxQ9rUEck/kqo630+QDF
PKW2bG70qcE5pDRwp/UJanfeVqjumiGxth9tx41diZmoEu/2+UxfCQRg18XG8M4j57EIpjyQY7OM
1tYWhic/zVUSbVR5rczwGzPYc6CsR5uH+Hut5eTGlW1LE9EwY87xW5VnW/MsOyDmsq+gRZQA4pPt
/8fhvL6eIRnluxhpgwTVfOZnGZyLqJMOzTj/X+P36MaAQDUP5DtccTfPaKXKXMOSVIscjPtX/PkC
xEf7SPbNV1Hwp7mnOwnUgnP1yG7BDF4BZLBUR59qvigCwO5MLS7jbZvfZfLGONmPlMyCoBCoHvzm
zEaJiXYoHW8avAhSKRTVunRFfJ+D6JXG81OeyKXdArtLxSqWFsH8L/eOiAJPFXazXOdndOrhFLkv
CaSlZ2GODzU4mdSmbGovYwVzAj8zcseP1DpmOoZ3K3NRcYdm2pYVN4SgKrJ6OwVsKaIP9RWyLTD7
v4wHeg311WER08wdRGqyJNf/QfcqPV6QoGBSecnYjh3+vY1EDPie14BNtwZ6tREo2AM4x4edXeAn
qhL132h610+vj2a8Ys8DM8T/ycySV3TuhQwwaNLAAIGj1rni81WCh8Dj6AniiQzc9a/75kJbe4er
y46OsXnVHJF8j1ykP9MYZmwuwVwIQsPNpmczWZ7Asriat61G/0pah2wHNIsV6/Wj5ryaKZVqrbEc
gQ1EuqHDxzeE4Xhk0yMhUKoY+qxF1oJ/wtoPNBkg/DUcvWwwBQ2IkhWkLGEfBfATqg8LKKybWq05
a+EJKdWImumz3A02yxDX64pyhifL5PC8w6IFSxjcnIJcc48R2UDaubIhTEMobPkjnxDFmiPPzJdQ
rBbzJ9DSRpHZkxAkuVSy8o+M6mI0r7WEKJG8dhp1ftcZJICI56Mxxr1h6v9F7K6hlOq8XQlhVaec
YHJxhbk4xJflWOQ9ukkKxs28TqUihPXFM/vf1t82sSxf/eNCmN6ug2xnrsaaFa6dMGRn2Vzw0MA3
hsiL7nct/kLDQS3Yp/X3SCW+GbvqTUiLJTJW9jmXo3pjq415p4Lq5fgC5O/FWwCJVmhtEdmU6qNj
0y0/ru1iKWHqbz8pqQmY7P27WxBT2UYl9z+/hersB1u2fdd3uqnOk6nh0cs9tPqVJYqp+aU2XLJ9
5jhxGLSBepdpG7UTsyyV9B+x4FW7IgFJ2JfGedB3JEjx4DdV08Z/7wOJBd9H3SxW71KujOB/ln2l
G3bDW8BUQSiy9ab28fa+YpRqxUXkVpRcjm379qJCeprfAJHH3v3tfCQ3iaF+hNeZwXvKndVy70g2
y3Xjaimbd4QzCi3FTIZjn3sweM3uo9g2RgtK/Ybk9ElgRDW872blznhQPA+sht+s8MM7XqNRWL6i
3fgZkywauOEzo23D6wCECca1YlglU4dmuGni2NEzpMPCI10RfqToskkckYJHuf4MbQJF5KuNxl25
+BOXFr4HL4JMsjGUv3zU/3pB30Ei+B1Z0LTwshB1rgS8+vz41ScxDrLNkh78qAj5oQfhGU0w+Aun
CfQ8gn2v4r3GpODtIFRuai5DLb8a+dOOvIke4d60C8hJFm1Z42PaEwkqwP6VVeaZFtFwf8P8Ddq6
SRaIlk3Z/7r44zx7gphamlWrNWj3OhawNyEvjnY8qp6dORqshMzNDWSoDIeqDQHWSZtB1cuSGoWQ
2/s0Kv26+QWaOW4z26SXLjRIoEIRRmx2bMiorJSrEM98rXjuxPwfgju0Hw6ggR6+4KbnMzHUc5dy
CG8VqczPF9PIw4Ni0vtl2Rw2c0yyDpW3g/n/lCJ915d3/biZSvXqMgQHXlaUv9jvCte0JAhAUf3i
H1Hwv2jofwcg3Uhl3kkGPBzM8fpkKrGJYr3MrUn31FaWWVJ1fCjcTAHmLXvrRvOX+DGLsCibo1H+
Kp8PGj2Ma7dYckwnGykGxU/nIcl8RlaDEoDvlLXgPaAAneACXHp8XBMV71OsmLglhj9pL54J1/V3
Lv30wS5uMs/Q8rjudcnt0ucqgUPFqmcxslbVchh6UQcCKS7opxxqGf0PQop9/JLeg2Qx8oJ6d0BW
ELJVltNUeMZCpIJvE6TfAfMLShUczpl58B2PvF77ku25xup3L6hZR3hm1osc6TK+FnRC2/d6ZDbJ
CkCDzg6AEC7SYQRTfr0jcCQn70uMcOPH5KUyaTf/fY/X/ucWCm4jW1Hm29nP8XCouMU1KwfEYA1v
uyhd9z1pnGgFtKmQfxOL5XGj6drkVTVWjRmN2Jjo6VQbPlr3HykzCpCpJdirMhP7+IHTkirRztlT
ZfNgn5ZaiM2ncdzQ4cXGOyNCTp3Ejp81mJHobO4hY6+KKamLOrwxMJKACgNSC+jF7GZ9W9kz1FxP
8zHKWbStJqzqojPSsNUYbXNMpwuukpJncaRkIbf3N64E1tLmjZrw46OCT5eQxlhnWEVAsr8GxBPn
84/OusKKKSRRKQlDfMEDk4kYfBCyZJqqO5gUE5HQbAnb3kwJMeFmLSd51NRqAR32f5E/wxVIsrOn
XzODMuX7XdE/0rG0MkS88ubs7pJ5EQ/nR5KZfQV8D3v3ffVjty6zdipVc4S2kfI0CpgMM0Yyx7n9
evAPfX1l4wtI76C9u+6mlJ1mFfhHTYy3dvjaXxX2qxtYTD5fv0vrFzgMPbEKZR/UywRuCeO9YjkE
nG1AnD4UoEWoMyycjZ4BsiackfP3lAckWFgXJxmiqnaT/VSnRDyUWGyIKgvswmqlJcF6viSZa0R1
6u3wi4oGPfzwtO1oENeOV+kN4LJcmUrzYE/sDTkN3FwcTPMky6if21YSNyryaU+W4jU2RbOZJjd8
T2wWNpMSzOmskqB0t5Pgr7ygm4YcqTtpGTY3w25/Dg5PtwtPG/7Xf+n1NF5GOVwjni4cnfRQ0pY+
lYDw2UVj35TCN2ocaXwFkEnMPJIjA2MyDiwOVN5P5+/nPMlx8eiZwhyalTg4C9BudW0wwrN7wrKf
uFWVRAkWjjaE3WpR1DIVhxPwE1l6TMhIoXwRQogqr+D+MuUA6Z1CY5unNGOnVDaPZuFv1au/jWRs
euojgAXxyzONtL+GGaui/DtMH1hkU2HRBY7lAJvtlfKyhUdtVXJj5v/WNqaLEAy8rtxDuv5O3lHI
7nDrKphxSz9omIvyaFD6KP2qmrfOnMxJSzPMbgTiSPR9UFtDm/tIjb8XMEzKy69yC1Xdqer8V7GX
HFoWivOj7K1u3IWZSFLpaAjSCUs68xVE0PWTFgx3tnn2AWZGABnLaUnA+5kcsabgTZLsUrXVts1R
Ofm7EUSjD7v+fQJwTGTpecrykqOQ5YwxIanL9Zv4tCu6YjhUEbPZzQeE0zkRIWXgyvPcV618bkiB
jlXHy9fPakrOUn2mGN3m+bFGP9Nn72WnWzyHkUpQzKjxKWaFECYYT/wfOlAG5ptHnFLtjhhCaKOl
OXnIE5R2Ngtm7o7oWXjoJ1Dbdl+b7NrEV3CyfslxJJjXD7IzOjTLVeFv4AqCoKshIBrQY/IYGzjt
5teuejSFH0XN2nhk9FS9TOZnlJqsRLls/ITmfoQq8P7Dh+9iqJZhxjlFI+YGwh/pCyodm3mTd4SU
+80l9CmzNIbc8AZeoID0Ntvp3aPl+KAPM+foU7oqhNvTchb072BCoLjI1CZXpfdUb63kH1wMov3d
xBl1JLphKEuXg5FuRqopa30BZZASgM1WiiJ3/Oks+w82Lo8FwpFG0B4yWka61q/telwlQIOUl97O
i+IHFQ6SS14lK7KquEWA1XH32jsH33CPXjSfi6uz4x/DQ9vp7yBq6hY+qacU4APPNqNDXdsw/faK
vr1FP860W7j6ni0beMFP4kjwJonZFfN6F1eP10QTZqfuAh8pDW0G2hAP/GLivronDiS2anWjD6/x
b2ZpOcr6QEzh94LcRhrzwMKZXmvQarKxADBb+Wpz/Yx1cBaQ5BF1zD/8RYGJxsO+H6m1cuD0R9Vu
qs/Lw1p6A1Td0gOV8GCONzYNftYE8KkxsYvTY0LaszKr+hmUY0XPi6x/Cbr4R3wXHrHFvHAMEt73
KcwY3IjZIG6OsylAHUuEcgQGSBIAhXmOUaN97rCPQJGKPZObmEw6I/RagGDU65Bq4iKfdZPDrv8h
VgIxCsyNaSbm23r+7Y9nortjk3qZ3Fen3tVar25Esv4Bnww3TQuXEPXfHxfSaQI8LRBk0xb11WZK
2Vj0X+9xr8ZB0hqWiQ7rhbFNDg5EopTjzGWuimQg6C9Hr1ojVBEERZhl+eztkYaVSn0LUFtiWO9q
AMUJhqksAFyERkQGiQ+1lDGFGwwtdHlzEyoH4OYakx7Do/nfji1qX0DU75tdOihULmosR3kSYCgM
rTgn+/EXtwMjNkS+sH0g320UZQBVkJoWIitDr+pYbnyQstD6RaYWlqlGguRR4KyhCrPnpzbYd0U5
1Pf19Y1uZ4/dwp2JULKLSjYwOaHnuNZvue6X50eeZG5XWHrnjYUPYcamWkqpoM7pGOXIWsYEuopc
MnG4Qm5iNlfhfOae5WOgTTAtLux6rEyUSsOReCRd19P5+YwwhgWBsSQUXsMC2JagbOD6ZDl4njmw
GQnYbGhqlQgrqWPwatYDD+hICZ0VFmBC5YyIl9Jb4+OrRD5t+JV0y2QjOhfe8DUG5PeezZNLF3EQ
0CErx9Isehl7Fk+E/euMuwwsV6SEWdnpLQqO3NjLJ1LUWT4RSZqqNHsYR7b9vNoOOviCvQ1FYLFP
XmWR87f6ylipJBSKmbcMYqGpGpxVz9pp/RwTTRF7EF/DWFYNnqAuOE1VlhzVuIuI13f8ee7+1Kvl
64cbrV2GWiZH/iO55zjOQM8x6VCoTpMEhTks8tETBxjMlKOlb+fGyCNu+8ckRXqh7QuzsKlggYR5
zx94DnDCLlDc2UyuMWTJlU2cbvG8O8beVg03KzLHFkD12glQnot4C4VE9XQQHxK/asLu/aZLX1Xg
AfG2P+wMtlb4V2Xs4UBvY/VImWm3kMB86zHkUiA6J3uqgpAu07Rfs9V1yZLeZiyvLXyt6gFitYVf
Mu3SnylGgixm/ECbDrimJKi2dGQbLp0ZZCQVSpEBL9MJ/yYvEzrH0L5D9tH5Z7+upc5ZlQCkG+vs
PCfZTUsWlrLu4SmSLzYuvd2XWCNgOjx+RAmtRB+4P9hdEshIsq32MgiE/4Oq5bwwywkY4bpf/cVK
WG7uPdyWzJaR1X4jJQmIhB22DlNZqqJ+NWK4FiP7GZvolFLyJdwQTh6zkRbT2WVTDs3w2AW06oOf
vAcLk1ShXPLuAJiKa+h68Xbuy+KpgI1l5UCpCMMHGfxsohdvHezjcLNa7810HWg2QtLutPnH91pu
SmLyuKt6AfSMvyFL/xuO5loFBwTPApCNLRq1wHpLlui9YeeBhmaAX1jwF6dNDkRPzlurVsDhLcQC
gjd0uFTd6Ek6npFptRnkWTnwuw50dz/6DI79nWprdcJwTweYsuDcj6J0mCUa6nYBATcoecBlKYAx
SMIKqwYIw2F97JZIGbdi+/gVXSgdxsFIzlrgoN1JCC4aOQ295fc2txsE/m6+jazaP7MVGp2KoXmn
DgmfkBozeZv4ayqSnM77AEkXptXAK9+Xq6AWyE/Q4xN0ZSWwvfqYzBU5evP2lx09SmNJayOErpgX
1GeEHow6fpAyRvcjWpAW821qzR95NwTrKEjDr0v3YXXQ+kXMdpBxJjY1PKX6TwkQAqQZw8Fju47L
cIqetEUS0AiPb6om07JPn5I8UpCaxP6nYHV/qNYApBUSjU7BRKM6wEbFzUMT85KqKYwUsTtaQPXf
NNZRte4LWyjbrhVk4G2UQozmCveghA9h6isdAxhHTlN1KZEFB54ePcueW2mtn15wltrGlO9mjK24
KnERrWwbaFZ4tfYMhGl8Z581fy0t43M5WTtlqq/o7WxMh1j6g5xlF/T6SNktRwAfN+W8NaCYm5lR
oyQtqcbVBCtDvjiC9GTMS4TG5Q+y2py4Q6k+AcKPT/ZNavSMBFF6Clz6qfUmVtkQK0vhtTnDcsUa
nZD0jn4uQM4XIB6hK7NntaljGcbjfAKWR1jWYkUapPA/n1ZqUEo2HuUniNX5awCrALsI1dgpLV1/
sImexrpZeuLFcxbK3IOhUKKYfvHNkytj1H+yqyJa19cI4xco6M3+BJHhM8syYXb9BFglq9Hn0OG7
ReFae/6gnSLxZQazRqXLVQB5abXm1WB+AFgPjVoTjo/yk0MD7vkBMEqA7czMmgbA/nFrZTYcl142
HNkCVWbESkMQVx1jrO4lvjrOodSae0hzEeJiCmf7rKcikhcU+0S9e31+Kp0quPgz/AhgA1Plufbk
1iSaEc6VY9zr/TfORtE/IXyra2ZXszOsGr5SbK4mBYcjTDZRcKffIWopRqMd7ehVDcH+x2oPUq2b
YQm55r3gsE6czUmWp6W/EMvznSAhRLvX3U8QJ70ksCeXOx4TWuwQaulPIT/2FuSDtxj5HmWp5CUD
c5Hdb04SppSAwv7X3YzXyJLBkUfNCpJHfK1yxbI8SR1H3t56wJQBYk0kezSitnyPoW63yN8cXffi
7+90EGI9DvnJihqAH9PK6E0O6I04+iQo2wKtLOToVjeFXdg+aPRTaI4IhLI8zSICFgVUPlybC5g5
EWcbQa9baR0ySN7o9F1XQv+K66sKuUjlTz7eRu2V6olQ9omKoCKM1NUXQQY9JPxL+az9O/TtC9A3
pWD4cEPpQ7W1/sxPkPV8h/tXS64aj70SECqn4r62IM5nUZ9jDP9f/IOfjFzKIP+Vvb1rgr1pClgf
41l1m+N6xnLiQQmgA8ggcXbksOIHqImq2t0eUvRFj4OtsIszAkOuyvigUb/Vs6mKNWe2d5vrzF/3
vHNA2Zd8P7z6SZyZg49YeeeTeU4Lx3DOO/HczkHNoJGhYZSWXXMbZNZywLS+infiEXiZZa3QAY+x
qQkidfHvVZD/zCmDsCyqLuarAfg5z/ENCFfdUB9TG24LTuVKUJuO9hRE+EVLy07x6RgI1vTOw88g
O2JZNAu2Bn8wjhA1UbuyE3i5oYB1qjpXvp8AjJBytrem1ZfnRZeBFKFDfePtk59aAz5DoJfV+4xP
SsAzrN0AyEFaWcvh/DPCTEQDqwkhYg3FMMjIjJGflqvwqft9wwgZDAMGOZdUhpJ4EJ0fWr9zQ/DB
WtZ4fHjCvdnh1mm3LQfrVnGhm7re0K+Hq/Leo35WWo+QZe82pcRrwwA1JZ6n2QUM66TvLGnQgN+l
GZSo1do2YNWOx33QCSMTi8FsUslKDq0ns0ma13ITSeYUG3Ns4mNIYxNgzH+FeLwV5dwnun5/b9Rp
wTIevTM2X3fWUhuPtHLA9sahN97LETabH7X+hMdBdm5iD0dB+pVIMWBH0i5JlSbBtB2dOoTNl1v1
FWdFMLjyXWL6Tk3F4XCj1AvUyaO02Xn67AOiv6EAPsrmL6svFH/0TPaHFraQ6EJjmop7Mo/bbCpA
lxCzEwG07B+B+PHeloBkNC8dJ5kwYwgeq7Jn2xkQJo+I7ATQciTXwSWAhkKvWbZqK3sTgXlNjQzF
lNo7nzG7x0Tqk8uwW5cS0l2/edv/0VNdxLKQwR1oPHa2dtBF2a/PYJXnSNvheWfMg1/2DjjrjrUB
QGPPHICgZhTJ0aj+40WqaVIVVmf3YyeD1bVbfR6ffDO4b5QiOmRJwYYhUQnZDcmaG5tPuyrDqBM3
tCJeWF4T4osmoS3dAO2D27fuJ3m9jPmeZGn0n9uKrU9AuIsXUe7KqXq8ydFlp8sPKJcLxen7+TI7
kGMMZaiYj5sCOr2xqsa+8Jkvzp5OqXKl4UmP92sAjiGy7rLISN0BJ86rnhIQnJfPiJoGD+To7tTJ
3Ya/ZYCgXe3TwWEwO0sDN6uIGNkslcodQQ2Z8QU5p21LfPLHoyXQeApg4hNrNcqcMdhduyynRaEy
BK6OBGc5xSLsVo+ExAGjb3Eq7z3Z5Eq++dWAS4D0EyHgQDBmjK9HpvmFjhoLSQCPnRw0I2A76ct0
XwsD7gPlBO7Sk+Vsa7SdeeqPf+23XoQDT8KwxsFJKZqUObdBL4JVvgvXvHXl95aPPpfuu92ysgHq
WPr4HOwObU0BhYWGxt6rSZvYhu30U07NQNLYTM9g3tltEWKNfxMgoqi+up2VNYCCNuRcp3PL2hbv
D541OgjfV+VSzIoUdqT+SmrSnNWnUhObdWj9feduhc1sAJQZkJtnnk49RtKf0EOWkFvsmWSbCT0T
y9HHaSBCwiMrNGsC4/u3rcbSYDYKAc95F8OPSbhKKXTG9X+2pXHhE3ZZS854a06BHpjDQKQWHKfW
4tIt8RBZvj6h8VYr7wJ1AibsKJ0qzlNhx3BdsjMktku8SewH+EPVKsfYatAwVKdO4U5uj6eIUTjR
5FtVjiSpxkBCQYC94qmjMXvviHWDi0s1XB8qYSZ2ruKUP2DEkh44iiO6xbAhUGkNWva2h7QIvRkl
pzwiDWETxbDIWfIl3xqAOtM1XLBpRqa6Vd2p7Ptce3VlhkQ+6isaJ0qV1OuC2xg55wpvxUUxwi+q
lf/491xt98AFzGH5WjUil1G69Ppa4S8D2eWkGcq6wJaUN0GLwD+BUnormXeRtNyqOBgnCr0Slp1Q
HpKuVSRCq01mjCziROJduNnMzJeny1OIOTWJAn+TAN9B38tEvH2HHHFdYOUVhGIUD0ec2eawgw1G
ejCQN8CkAY9ue/ByApwKEy5tTSK+6AZRiBdnQmf4hKM3YANILWppVTTRJWkzxMPuIsYpMSlYW9nz
mWNpN3zsY8dS7Y58w4Cxn6+cEvOw08neai0czxsA8owPwlWUEaGFkxEGisBT5hj9mVxoXhZEen7P
KPmxMUEsli/FiP5Fd03Ok8MhyyInWqx+9vziO9z1B0WjwadEZfT6Uf+s3VePgq54n/gW0/QeHzyl
B6T5QXRhU9bWEqOSSRnxgsZfnCbUk0aNqY7jDrJQStw8g1MoPV0wQ0jYoyUHkX/ivAtyJqj9B2Dk
Ycv3KRh2GMeLJ7d8ptEDr5kjtt5e6Qi9Zyzqf20TsV/9NaOuLJ+VrR0YE4m/yyTpyynXNGnMLAS8
06TjiAQbDF5gqUtvMnPZ7votjyCHJdRauCq1IrCGuU30mwi1jh/b3+OvzWTTZLqA+ab8aF7gjPSR
QtzDRQc8yldssJNndlrMw83+x6agviFwqVeKErFZc8jOyfzGa2A81u6Clpr3leb0vprt1d2I5ZIl
Lv2MMi1GUHtPNS06aTTGAzVRP5v5YuldZLeKBIH3fUieH4pOHBTpraz5v8HxTFipRQjKinNUWe3A
+YDAYdvFEadctkk1+WRH919OhJnU+sN6EdIHMYo95bScnwbqZ0CHx39YAFUZk4y0ZwqS2kokLHRl
gYJWo9hZQr7AF1RaVkp5XIXImbPRAj43VYfgwuNRlOJ0JrE7J2X9nWRMF4epXtW7Tw6ta3N6GYE2
jVfDjP/2k7z+cCwlq8Knn1uW4vQkPtUd0DxJqSzuNbpQFzeeBthOaL6MNqF0ewnm3zwzYTxpJgTb
pSB4bev4ffzBzsejqyAyH8VBR7swNL5SpqhL6BFzK2DW0kofAtp19nBxOcNQQwyaTF4Qk7jcnpoK
Nm7XWjyedd6br99ch30dLOfF8+Use/0saxGSd35H5Emdf9yFXrYFC6KxC0DXhybr9V1F4xAP6pVD
s+oYBTuYVxVz6bmMo+u2U6Vk24VNGb//ZylJXd33e4Z3okgoAHGY8caKQX360hpixoKg2tZdr5J6
EWYV4LA6kBo65aaMw612khAVhwQ/cB2k/lKe5VwFZdKhAo/bkjTiAReGkaxkWIq3nXSdbSXeTyjb
pLEcOsuc94q1AWeIr92WD67iQZVBtsQVO7+4q8sLDEO7fsKUMpgAY3Ho6KnoplXv9637JihPSE25
E2BOlw4rIJ+iYEd9zwtx87q8Z0DcqC7+hFaTEIkkMFlxgBY+GThlEged9N6YlCJszrIZ0KkV+8Nw
QC2lzOaW8AfF3GqlRajYgqE4Mc8XIRommJokz8a+NnY/S5ie1uq0VNbgDS7No2TQ0u3ZyS7B4A9N
GGzrNFA5NCOogr25tEIvY6DWK72CW5J2TkQmzc5M2hAaK81o9/QsVN6tti566p6QSiEWZpCZ0nnf
fbD3e/dZ7L0d+Pp5sOiLgqeaTNzVCElYWelBAimZtLbxvr+1xswHmiNof1xTNbrSThrPx+0HvncS
8cxrU39wI99u4q6ThwudMHmFSzruwhnmvb7J1ln6atHtK/fvtzZoMlxb5S9qYXBI9zdP5OxQolPc
p9Vgn2NzYHm2XouIJ35VGIajrL3ZesHOon15QAMkL/dkiMkMXrrl4VixiqlkOUgwW38ANDfZyfp4
ZWEL+ndAbo/Q+dlqtGLLJrnG0v7rC0uj3Dp+lNpurBu684C9On1bqsDcLAH1ia13ojIRG0C7w3Pw
AlReWiOzJOVRJAsP2aQSLVgMLUmTo2+NWtuvs1iijvfGr9VZgNgASOEZXls2UKkai7Qf1MRql0s9
ZSC/Uecve5nzab42bFP0TDbZQ7FNcP+7GRCX9l3pYNYKRyHnpvz8uMKeXp/3YAXllZSuWEsKO+EB
PxQtAtmndJk2FKRfP1SM8lcmZ46o/PUPG8LTFytAVItltq7Xpe88uPSyF3dyHpj7K8/gNGN4XeCh
yuGR6neFIOcnvef8d3Zd9O8PkG4wgPUgJnVkJHgTE8WY3bDbnTtMt7jLIh7ynfo9GHia361MlDdq
c0Q8nheKEooL46sMmYBGntavM9ivu46ytjlxguYI6P6hCuCFVxGavEFN8GYwXmGdfF3L/tckahp4
K0JwG7tPDdRa5S0dBNuKn9ZbARcTGb3UesgPcPBxLyCtCz3iaH2+Xr0ksxMMCJHQ942D+ZjInYOl
O6Wn3gWH3bJ4IXARU3qrxDCazN4IiAM1wE20P8sTH58gv7scrUbomNYycCMxxb0mslku45IH60Ms
UtdpNpEQnjgrOYw0zFSvbBE6oFmAqL+mYBdpuYRqDcFU5Q8GC6/GSafA8ybVkyDxZ0G5n4bLeuXT
g1YRKA7hVjMFMuI7aCkczHbcbSu4SCwwJlCqOyhs1RokZAUq1dXS6Yq428x9iTR0v8FXQj6mxbez
RAU5/w8JsGqxeFKVOvtaPWwWOjTXkDcWuMAtd9YeHQuMMlnzxPS9ODw3vfyZhkxyanHGS8FA8r6N
uvh6Gbds2m0HQc6k/mMDDs31eErg97ad7i9xJhYTQDvezfOVoXVx++GbO0v1a9rmWWRaJsgry9YY
O9MFpUywdDhuh/5f0oYPo5mm3hPlKrmFoefNprLxDth+IuTUQTxEALIISMnsPyrOU6U34w3J49gO
kuR+Ikjmz4GUaM00vWr6U1H/95LHjXK0ZKzgDQpsfMYd0Sg4LGLP6nMY1T8Eur63fUoCexgOpELK
SYCEMYHQnfN+Kvu2e9apakQHJLTyu7fq5pMTL4qE14EGFcZfWDJNE5Rz6DX7naiBUjFSRnrISxYQ
aj5+IzZGq5kSrpk4C+GVJLObPvZi9PjuE71ey0Srk683opfGBQVY7kNPTw5btRpQ54IqGICmQ5Jt
mbtJHDIP5FnGBIUhFQ5AZpuDmETvhLtU0jjLE80/Oq15SNss7RQ7RIAgbXsCDa5q1hoxlasRvwmj
7/jRus4N9XABGMTUEfKfsRC25ChbtGJIE/QN3/cOiACRkXXyZ0dM7Pv1bQVZ2lLxQD30/vGi8caY
ki88T/6XKl4z/1TcufdhbqvYfKs0jtLZQfHvZbT5Xht1Fdk7pnnTbifAWhTwD729sUncr4APngKz
ZXtRUkAyfj0Uls0jcx+V4kzOiqVtbPpRhgJmpPAH41oq8Z9oE+iaEBwhalVKpQ312axmxDCf6Xnw
gxqUe5nhonH9xh/6m5oR4Gl8bjYL9MkBXIpk/EdQmzOvV1DdiaAqNf5lOwaDdHnCEEuG7V85keW2
WuLKV1E+UemlAM57973SBn9HlCgeNh/WEB+kfbMguL/3Jc/+ok1q+LZ4gty/itE7RomET4WU7awc
08HMvbLDnrzFU/d7Es8twfPEu+Bel9d589ATNFmZpU2FvOytWGGLnv9diOLRuzjLFnXLt9jyMjWZ
PHdPhLYxj0oDXsMR4svv6Lk5vV5/zJqI+gJhOIjk5txFENsCJD3XAaeNZeZ7p7ENCVmmFb8f7G9F
EaqijAck+2A8Hf9jAYjK5RiwmjpVa7Tx6UPS7+ZGbelYxSik8Lsay0fHHSNXrBgCE4ByfNX8LK9v
w/7/yWgHhuWKhtbFoqpwmJzmAeP4UWwf1o0yIabbVMYPIvcLPGoFHn5x4eIVh2SBbxq0tzxyHlob
DWqFiq2gjRQGvD7qEVRBb50NzJH6hZHKEjOgi4/nwwVJF+e00vapgpzM3hMcuvSWhB10dsuVFOCh
/7UOqExWsvPQ9fN/WS9U1f3rTEqAzVnWmehEAbTXkNeitou3tdCa0EAIpel86m9Rt43ifhEtvMfa
gsh+EVtgrVAIi4j5A6q8N/T+FwH8Fky3dpOL5EaL/UUZ4JZMhTW4SJ12Z0CJd+tgcKE1hoquYEl4
UqtusOLOYVsYJCK+9pL6VYAVMCuFjrbl5xiDcuUT8n/zIgTKpzZkVeYtBEjsjFSh/3eTIEzcaQem
Rkblag6zl4AHzOdd9KPVL2DDMeRena0fzUBhUHEiihcrYc7rN60vEUVBg2C+UMG8wXANMr5bVaKE
2EcjoUSJRtil4GzKrFLVSm6WzuhNo1GgHpaF3tZbylzA9CIxoNjsfpEaB2kBBRtPRSaYzzggact6
CBrRfZf7hDjdWfY8CWGfMj99P4VM+WhD3MGtO0aD3fvO21py++YDZSj3aJvK3eU1tpg77hT72i0z
MQlGGLoN6Wd9z2FV+IZCuVP5EXhCPBph4jyDyXgvJsCyQ0P0VCqSnCWYNaKTqUdeo1tiIXnWEQqO
GOwxAeti3NjJWPsSZs8mH30UKdAwnhkbNvCf5pZ+u1CPsWZsvGVhToG56KH+nJGjyisebzN4PP8/
pF6DSCWTZQczCCjzuQ7hEbYWgo26G1K5N9jfvDY0859tTGXGAnTw3vP+NXpPUhoxtrXRjFlPjj7l
tnfPi25STo+rZCkBVfr/+SbShtmxdi63xksguyLrtmMBr/Vkjb0ue2suJZgHw+ByG1FlaBq/nUR3
UqR8LFi8L2+PifilTWphKKrm2BITWZc1Cl9b0bUUCiLolMoepVw6/szWULT43+dAiUvOiYERmWLZ
rQi6UJJg4kyxP7CoaD58bmxTr1HIM0z2FKau0HPPlxmYyXe+vJ6/aKmEF/f4veSZTdo6tn/f6zTw
jD6Xd0yF+537c8rdGrhllombFZpAScAzdWUfp7+4LlYECus01fay4QY4SNCVbcwuNQGvcIwvKT7v
fDUKz2okurU36HRH4wRXXyQ89aNd6SV6pP4AoECcIvjWeb5g8GkRdxFn8c8fMkTU9q/V9Zc/FaTG
Le4wCunHlQqyXf4IxbAthYjMoQoM3THZDswu8bkBybVc6x3M3RQo/XV1efQwDzanijCif5Wp5ZpP
OJcljbFdDyJlM/iOe25K8s9mywiK1N6qLMmJJmlEzi8ej+RpZ0rbE6bz22MGKH/fYnCRvhKV1joo
xAN0GWu6ML8EFIXixJ/P2mem7vL6NY5f2OaiMXQfS3VLPNnNsZiPpJcigw76NwXKo6//R+yMoiPS
wCv61tuhGRXohZjhAvsRl3nYTHBYTQPNCjLqpV71oHyNWdibIqZw4j4BkuB3GaeHDHGHpzUt0KFM
F+mJ7jZmZY9zNaa8gTwUmCXqWulo9Yid7DDO3fPbRq8WX5A+50eq64zPUBOvgNPG7sHb+4Y/743R
BkYcpmTV9Zry4aITIbpZlbKOKNRZ+8CGv6iYH2EQm69vVil8wd2TCjkcP2gAj58d69ZtB4QUmAXM
IXKlx6gJgqjExgwMx7bFO1CaBLvmyA1owfAaFDnImxLKPQHcpnuu++/g8cx+PBntLNq4eBCs9eRu
2GOGXwYaZqREQpyrCEpdavfbNMequiIaowHxmuGSgxXOoz7v68FJ+tIOAgoI/FboArz4qUcp6IRq
IXvJSkRAh4a6el6Q6zZETJfIuppcejE+JeJJy/0mzXoozdpVv8NtAEopf9LA1ov+RKZLqG5PTudp
bu9dpbd0ICndUNT5DNesgr7fepFNaHly5ou8wI949pMVojVLb6gqglEClFXi4wVPLgOdh4essAhb
YvqRKVfjCVavfT/w1FnyEEdZbSL3sK5FnhDTu6auBY1HzPQtkZ5ubqqNFklLPDt4aRcV1O7UXGkK
5c4MbGS6A1yrvJX2fMy8jT8I9gaHI0uujPCUfeiUgFltZ/vkmgJE+0kfhQ3YXyyJv8cM13rCGpJt
uqNxUMoMnmcDbO/NYxd1TjZ1Xxn97o1b68OcoJ0wMz6nAN7Vo54owPRMav1ToeWRFEsWUFnStinq
/UfiVyyh/qY/pv5J/8wE8FqDbI1tU9A/diNA7RPNPiMjbdRgnuG+pMGYTNGyK5LrVGFcP2d12qh1
zT7Men7+WUoihcgKEKIyJwAt5kSOMlrsvLDdJSDS0WQuVUOGKs7SPwYtYAcqxuF/7aIjCyx/uePu
a4YhYZ07cLSPcr5oA9sa8UgJOva5wkQfOHesKPrQnNpIfI4AT9WehM8inwx8AReVFgcyA2p4HeLX
H/rCCB45atlINZChH8/tQ7ZUWfDZF1qWG0mdnyvR14OSHNVBJtMXYbGIVR7xvAVDXjUASSjMfDqP
ZYfU621KUuyHgA0w+gbXvPJohu99gq9AosMtvTNzJb/dfNVhh6rp1WQ9FwfKgxttZVS7V2QJLkWF
jQ+MwDPKF9Z1BkUuAe4UlZijp0/b41/2JY8dSGklAThIA1yCFNmC1jg/Rut6SgIwdkxebOqF1bRY
wjiGtDSDl7TPnIHuupq/CTV+E29uBqXgeUB2O9KH3obaCxcKJ9aRlk9D2bOQgEaG7vQClJb1Z1BO
BKON9DCo1+jrFcQdaFnkdNPctcICgiDibbT9+620HDudm8OpsiLcD+WHJB3ubydisA1H2Hxk0sFc
2p0/g/0lVde/PxBaSz3zaoenVuNAbE/xuQlVpPGZGZBpF91vmQx3BnuvdwFd1YUAIk9yJBVbVjg9
Ce4rxp+g0/NRoZzAEEBcAuSJsog66Js1uDkHie++4Du9fixDIml7WuJlwtTPz8oUQeGXRcjqeFuR
w6vb/jdjEBuDChdUdZcehbxdeTesv+34v6rhvHCBrmjJqH5ulQbtYPpuJ8ijAQcD468NcQFyJu8p
/SsDLrAAXveXSOTuZgzwgOk8RvHmFWSUz5uQVRn3siwbnInZ5oXXdkzVR4wRSAOMqb1GOKWtHHYo
hx1iCNOhq9y5ZE/Xqq21gA+VgmAd6YjTRKbCMpmywJyPVtaUJqCaANLKwLxqJklFmVPxhOdxAYfY
dbg+iZy06E1F7vLNPYAFTEbHbDimgdDlDgEpV4DwYzcejOoeFe2GVb/OQARwyV3af7VgtX3bKSNF
/25fLZWCiG3O1ze5arcYTHXYwy2Me7zZj5h4vFg2XlkouRFQtVKac9L+yv6MaqaYltbDBe1G8aYR
VKxk/iJpbWM85MqA/VeCV3XfPmW1hwxw0xzNA3kLdND6XWP1EJ5krzzVk/tfb7nFesyPyLAH8U1a
iUYua4XffZuGyTvkCMrzc1BzkBdtu1kWAiaD5dOSHWDK5kVKWCAHseBIlKtwiLoKa3Pq0WT7zBzo
IuTXbZRdI1kJ24O1g7Hh2o4q8IePC4YkwWwi2znYn05BTuZC27+0V4eswO9gJMsbq134W0fsoPmI
kM8Xw/ZXIXrQPWbDVT/BPB60+Dv3vjWvWzMZP0bhaLsQvG2QoqQeHh2KcznQ2TmapclLO7hqRFrS
mWmP5FP/gs5+Rx6Rh62J7VkJiczXF/9y91pUTfDcd6WXYp6+skGuZa/gpDN/MWRPZBzUGigYyru5
aXrhypXC95hJjVKMWqJYij33w534ujfKW2v5RGp6F1MQWzXsbRlH2FxnMZiWgnzCTux87oKKubUw
Vjul7wqjKBOpYHmTdeNBV6cryQoXJ1wsSEMBJnlmvy66UXQUXgDckr9DP4VuEC6H4omOQ+s7Huqi
9GIIwmlzdtKkAFo24SW6iknvlNdQhmT+9vVSW0q02LbTwWkcxdPK1vQDnI37hZwX5BpX8WgEMUd/
Hm5rpbtsATNfx2BCB2o+UGCkRqCD6tMkybR/ro1aNLfSaZdMi58QQC3wrQ3ITs2Z56dAb+g5QLnO
RtiPvsQ0nIeJqSOhBeOCsthUKB9XSBEGAUvMs0UUxJFqMzIuPH3yEgAWUK4V6MU1gLVAARMxfvzK
3ClhpziC0FbuM+ikE4hF/ROWmUHb1MmlaVneq9MtgP/iYK0FbCKa808zbJ/Z64UY+xzdSQdZcHtj
/POEmFgRAkWLQXiXcN0zSnk/NqHtZQiP4KEJ2O9ruLBEPn2Eue24unfSy4HPKhe0M4OZhbFxdHyN
53yvlH7terimmVH8pKVdPjEjhrB6H2huDqbctuiCDJGJ12JAdQSSFISPD0Rhl5hJQUbqwJO1zeQW
a7Dd6liCEi907S4WtW6ehDL75wzNYmgXu+VKBPGdPl4YMLEPKHGHahmlHUIWfwa0le6Hfr1zT+rP
NRLBCE2Q0MZyuOI/mw4To2j9xD5PCI1PXW0r+YkCBubuSAwkbGH0lcwN/qp2ct/30yZJ1tujKren
WziDI33XAo3sTtcBKDShdVBYr5SpdcEFHRy356ewE0WBIj863xJMoIps2gEzbvbuliLXT8gAewMN
mdEpvVpAin2kMvAHUhBrdDsGJ7e7dessZn0SyZSzcMaw6ed9mKorhK5Cdz+tIC5tUs1ObTZnfo8C
rEVB6slVXQ1upq0w3Zb4z3lJtMX6y6AMutPnfDnOR59A4J6gueeW9G8tW/XPhxI+rJY1sm5D4/RF
gN9K71CKNmmORr4h0QuMrJdrYtvXHE2XhhC+VTpBRV15/pNDszw5XRxeQz1tsyMM0rBsxzLSctWP
SoDs3Zcmp+mOolu9XiPISu5eP9s+0TxABah3qPUgxAdN9tdfTGvzyawZJk67ztb0CvQaBoxy/m+J
7aQNJhL4JVod3275SOvdZl4Ha8AjM/znQBLv7eiyG+LkYtJ/mOOccqPW72AHoIBry2OwXnbhRGY0
BjOQ7jC9MvpyrD0wvkm3dziwrJTqvwr2T7rkNeuBBtGc1gZpJ88ZyrmAbKswV1esdZ7b3HVfFeYu
Y8IaoQhXWwJF0yHkR6avBOJI9YiMd2tl2F9e2nrkYrYO4WRz5OyMfx2oVNtdI7bLe9JFGLWALyPT
ettu1ZIXSWkZH8ND+STT+HRXoJ2fBRQOIjxO7Q7Ern9DPSexQ5MV0JYwJmfKjGh62pcfi4CFea9G
72wwGuyTIA/J02E/oVjJ8FtrXVFFJmFD3lQkRS1Jc4reJfGb8ahOM08UalSEcFbmaqKosQnZlOVz
RW7SCvTQr6BuDBHbazRlum2g23/LWeSpw4C2fQwb8wksUp9kVENj+Z5tqGIwEjBcqMb1ZESzwMnn
UrZoFdyfORzM2a3CH1zqVY6GUASu//62gxQcE88xjvLpoA54Km78MerMmlXA1L0it8XJXqgd0Ib8
vK43xuMi5uilNNaopZIjkkxEEJzamkuypgZesDtCDUCv0Zcr2LBwU3VNWgbv8yohml1Hr0CqjS8R
2OO6htfgpPDWSTVvchmlxVT3jpX/CDztheY6pnXmiJXwwim/2vNTdVcSzcOVKTY9P+0VY13YNldG
in4KfTCegaFHNOi+Xzygv6yWkHFD5itufyv0AGE+RMWXmaKbbc2tflXHmVUFQfwfv/qUyjKkxdLY
Ll1VQKKjvJpYged6QCS7SEnSu69Qd0rmhMDJzx2eGS7Hfa5Jfcfp54ksiINKnNjzl6qNCkbj4mT/
9D77ylHriFbf5LyToUch1OymxyNZptI/wze4ADAojqh+hi1j8689Ufa96OQZSbBKtGNfYwWEyPb5
u9CJeSjxAE/ArKC38fqmmkGD4ZVo8ErPdBOjVev2deOPiJiYW7GI0aXe58pZdQseyqp4enXsl5Pa
mR6c3+Y2qAERt/TyWeGY3plEzO1Qn9bGvMA6TcWicHmUGIw9j3YSexM2I4meCdNEZcsEpIR4oulW
Zxa7WbB+x8c4qlWwvQtFKIjbGBoFyxI6lks61/UAP4eybTtsNtz8xmZ6Kcwr+5ENfiGptHmVagpQ
eRL+TO7KpmT9WxN3qQlGPKwYNdAqaeG8OXknM8U+acVZ6LTc/CdZWCepa/ljtpmPYRv15L/eB5ER
0X33fvdL+wiYwAMh4H/EuEvgbJ5CO6U8WRTHifOc1WFVeRyONao+3AR128ZFDt1AY+Hrg7dETDfI
u1nF4sOCxB+aj3Ct5MXNbzYX7xVX4C2i1jVipV3iCxCnBelNuFxtQiYdg3uu7/i7gVrpDW2utgRj
9efuGKtODXVFH0NXE6Li2O3VqFumaaQikOqIfg0myQ37MfW+3Ub8dnWtkh9dK3gg0a95PPv817WB
foDHrb1p/ge62HA6unAH2YZwhWlW/VrUV5xqg50IiBj3t+uzWPIsvJRNE1GnOaOqL6W5fEU9iiEF
TgPYAfWSbw6KOCqQ4L6GGshMrv/FRQsgOeTshKCC4VBDtmLc0K7odQe4V/FzvmvHdp4+vMCVDQb2
X9zZ7dYmLIs5UBts1yMIeNVXSk82w7oJHcDeog205ILh6kVYq73dN5u5QM4PuikVqE0WiDumUjZA
4joFZC2/M5YDzIy1o3VvvWZjP/Huo1/IlSbjDroZKcpOuwphw+YUn0B4SYNk75RkDKeGzljvLWr2
aJFIRRQy65YYAFp9LmUPKVXEccg+/6KgeaKFhP+MeY9hMqELV/zUlAqT62ccjxcswksviJLi17WO
iE2SE5P61XgwewJwNpanHux9hWEPiizNhkX7q84rPajck2YryS19fKO58pdos0cbizRS7/QzSh+2
i/91tzGy4a8/8jaNIhd1mphM7OywqNICsEGvwtm5yvvuZewl8gw/nuY5xXGbtAjRebB5LL04GCHp
SD1xZC4b2IkdkfSmHdLfSwaeqiZjBnNzb1UQdNAlBjeeAdsqeLWXkSlJBLdB2DUAgEkFdGEK4UH8
LUUlqHCeoVH7bOabyZk1TP8kd+muzd4hrRUMDPnyPdcZgivj+zO0e5OVhsYVgZtgMMEhp/amNYT1
xpNdrWCac3YKoWHpM1vJGSRKbLZj1q84UGO5vQ/Tn5WpsVwE6l6veY9PNO8wYHaVa36ruH/LYrX/
YsZhIjPGzahkGnzsJw02Mu6rHg5d1QRtqZYKenR/1URGeOuDn2pdyw29efSPgwZ/KkbUEZDRkUW8
I6yK+iLuOjqQqsFLeQaRYHDZGVCLXUuXkDsaR6xR4TilegWdPm22DabdmGvV3VQ8gMN05iV+XotK
EHLst3KAvu2ZMpNFOGFWG9Egxi5hQWUYDLDKqXFLXccW2+748kapgNK+QRkUaeSdnByifX4L3Yxt
sDXfT/7z9Au+qWRwLAA4DMOa0t6jpE5EvGLOYic6aqKftrjT93PWSU6yAthtT7IKNNBXE76J07J7
+F0KBT/3QgW33k8sf/CLUCKsiwKeoDNAf+/AvzopRx8fSwayM8SjtMJggp6MeEWw6kMAcRdnQVpd
8MobuTJle5n+t5CTefHW//YOKh2pxkrIlz3Nex3Hxnyj1A/csdRN6nMpNfzSemHmYP+EUotI5/dt
QM1MHJDs2/LalGfQLw1q8VoepfGxf8xZ2LmXmwf/spb9nPMFb6EWfzGp05zA9rQyMHo4dQI1eHNT
vXhT0QfFSg3KiS/urog70EJ4T13vZWZK2l/xcew5LhzUGunMAX3iGbGFt6gsZEWiWrrpGaV4YK2W
0W0euu9QbeR14uNMSLaO6oCtMwJWAYEQVZOaqTtH6qHVEOAGYIxTU2WHE7/JU+yDypXUh6ikTop4
VhwRSVpj8fNwh3eUhmCa0ZpVlt3Z/7vlclrRR/G0zuFyD8T6r07cibB3SNR2wiJSK7l723KNPcWb
wGWFXOh4VMri5UZ37X1C+H2LaFIAaFc/EDWk3hL5+Nga2t0hrt+93nvnQTPKQcIhyE0oaSRWVwhA
3MbV+5LAas9h/Gr1qtL81Mni7WtcnohmMn6t3iem+OYbN7WZFHi5ZofT5EqC9EWTBgtrIec75+B7
eb6+GdQsAXW3Kal8uVLnMMgT68WwCLeEUsKM+9Jq+j17qp5tj6rLLfm/XOx+JAhv36wSNFe9tcpA
K+lYm8q61sxhM8zGyldfd6y6JW2KxGUL3W1XWNGoxdwAPSXOduRSDeIGssLME9v4Ec01Yzmb2a5x
8Si4v2CRa0O9Vzj/8qVXF+hu1fk8qX8ik9wThqEVMZpjRmGCSzDFUwCqvyJZDWAGTYHhbAD/RWBs
tx+EoP7MGgEl9QSws6qMedmD3+mF646RL+MNwvhuLbRQ687n44kSsxQBPTNunV21D3idQ8S+AVH9
lNv3H66lb8Bviv7Y/zVlBDENt2n7PFR5uIPKnwpIe2ddCjItuTrBgNBTQFvDudz1vqTT+VN652/J
au4txOAWfh8uAzWaEhcseH4q6cI2SCvtudNeM0/9ilnPa4GEj+9/5gJjm1btJ4MD1Ipr1JYEFLQI
mT3jQV7pu5YZYm0kJM77/hzf2m92VTnqTpi3AT+i9iVpKUNOwtbPI50lnm83pwk5IUZWb6/ixvon
RoqF4pvPUZxA4YPhvH9ZMdQJztSfs92YIfGkB16oFv6DWH0/96inU9roQXqvI1Qwl+Znq4i9orLJ
BtlB0u5egsIUT5kV7aX3IZJd5C75T2YhyQzcKsrfdp3e99UENWy56liJmTk7wZRd9SzmPA4215RG
T2ANuTqipWjYj9yXc92flRPCNMx6I0E9K5suNguPZzZsdldSV/yZnF6owi1lbL3mC+TR4JjXl7x0
6LaaijNahlJZU0aoP3lwmeMafHsreUN/frVOomTUcsGPMs5uw2TAhk4NYcOw/fLJos5uKFoebmwj
NldnRfh3Ai1ngxSJOcRw6uggrNPUDILe/07IbqepIdOhfIIpv2XuHiVqga34eVzcZHL2CQgr/qJt
qL2NU/tUXILSr3LVmH4p0ICnwxeA+vH3/fG53C++2/GjqOWqoTwu6W10N5BWnUsoDOdSzIquX9sd
J9WLHNeqH6FSwYPGFlRQYCvUtjy/Nj8ixdFEM4mwqnbwp9AXw4mLTQ5o0OhxeSFJFL9I7kqP36f/
bL9UzkVe57rIYJms6yHnLj5nQ+IOvFh4msBm4uy1JCQIx8pYr8Ik+g56Q+YylxVdbWc7l9z3GEIn
wLt+Z7MtkBuJHX4bcWuST+EIu1HM0+3VTLksviDjrMV4myzwjKdjDyvfn5wgqgTSj11KCU22NEF4
mGNNVuDQS759Wma82G3mbar+geMJahJrmIrkPxOyP0+lCMRJKSVX8ZtliRJVpHjGrYbfF4r87wL/
QIFDb5k974sHsVfgvW8dNjX24sH8LKQ7PPB1kiCu3mN6UIENHpbrSCCUh1CV1Oj9OJP2tgCXVJ1j
SiKIiBpyvDyKmc2/LnoO3xIsUHES7NC9jyRoR9SY1A0ntz8GKODFeeVvKGc/MollJjRMQfhHL+2g
VEj9CpnDBJ+Eg25CB3l8NQN1C0vWxhHrPnR6ELIRlG9tG8gg7xDcXSwVYwq6VxPPECL+nnNK/Rv9
/qkofXhBv1Tof+YuVIVJLElrI3J+HKpyFxpowPFUBVa1aX59c1mNvQq2M1amx4LIhr8Nj2M/Zxun
+ZvnaGtQqIwaZP8girOaFjTaSPAATFEd+kIiH14ljJPVC4XIuy2MHvtNO2uditX44Nu4BEpN9X4I
CbRW3AOl8YmpJD0uS1k/EjcJBUNmfLqKV/OamwAWHwPexaS0z1/mOD03g3ATS4jElg+DzwBbyZwL
YtcH3zluu8TgKR+vY1JZXmhLVDv5/3ZyyitzAqzPZID0V855nCmczL80IZJiio8xH2LB8j+hNw/b
D1DuqkDruM0Y69tRpNhFtxnzoD00mZJjYIg9pUiO1k6W2dcsG4doQlL6q62iSdCQU+/HcsJ3J2RK
Xsy17jqv559RQ3GKTdJzIR0XTKnbdIey8RuFvd4ld5IVtwh3OekyAMGzgD4B2vwAaqADgVsYEhmC
lXYiuMmaEDNdEkmf+k8oV6zCDdIh6EigdQ/X8b2fRrOOdlkjBabxNBWAHJu6nLnN4zpkl/2D5S59
rFvGhBEIsnSE/hEyxTcaUV/2wUIO5VluWiIQAuP8A3+17cMGFxsUIK02roq2xNG2eHzqeUoCCqXF
n36ACixcg3Lazed3VUIuph8SzrhC7iOtk8FZpgAMuFs19508ncjoXwcTFRwdZBSfZTAQYAu3XyVh
QD3P/3QHiaIIndZ9aL6STZs470M+Cax81+Wn1gAP2oI/N4fGNlMr4TfG4rA0toOQtHVuMUo1OneB
2bGB8+VRhsy83bLEebiNROoven8U1Qho4RCeeSEFjlQBa5/D2tU6jOY21SUzLETVMXdKgvGWC9AP
muwSVzUoHNWW1tVUuB9/Funv3WckEaJmJvnWXeTE5rORPMqyvlL9mVp7yEzdvzgurNe5/HaQV6fS
6jWYxqFkpmS0geIQmRtMi82tA6bSXY8UoAc6EmVy0s3yE0hmGcBgJ1j+N89PIRIGMw7mRGBWyiwl
pYluPDxHfqUTt609BwX9X3C29OjmWaJ8VjWHcSnGeW5hJQv1+R5kLlMiau9LQTDN3sEvsM/Ryvr2
VyNObEz9G0QGZFc5gTGj77Ds5/B0Uv245U9tzZ3RTIG6FtVaX3JgP2uoJE7Qb99/dZLcR8AdpjIL
dVsdHIViUSlJ4dfaL5rt7K2o5gT6RsZLHxr1qeTaxml1z5gTJPGnG6aU7M0GWSsDLDoob05/gMhk
jwjOUqGzm7x0rZm54PLLeySYglQGAYmn4g6LSGZl1JJtNZhXYo7iNgzK7ZldQBVysWQmMASPraou
ERDhIEipiwpBIr4ae4+fvQUMEgcUj2lKEDUpBur06B2+IA29w9pppjPsTosxO0i+yjXEh8LXdIaG
XxPX65th1Mo2R6Qs42XB/iMlRAAaFk/GUJzV0JyPoydwuXQlwqebvw9ggvVa6/PNJmG+EdiXznk4
dYgc9VHKCJuzLh6LFf9LQINeDx2xaBbCldkWxBE9WLu7Z/1hw2ks1zoS+2ZhxnAHMaV7NxrQEwGs
AGLO/7+xl6LnLcCpX4M6R41FMetdcT8sZsR7cG7kFbyuoSNhjo6Usi3oJAenzGuhA+3MrZ2Q39+O
hBCBSTsX4srVE9v5/VZxh/xoTjPiio+gdXCeZ0AUOgp91EFpHaYAK28hj6CFbskRrFpDwTgKm8xv
pon/Tv98rIKSrFCttNJsNn2OX3K7oUzOyUNP4YXrEv34iSBm3S9cNxngfsWGNEQV1zbMnhRN3LFw
ueSmW3UnaSF5ddscKCkt6/XoOjLb1d+3Fv5w0bQv1I8xjrOwv96NtOfZSWcwQ7dM5K1H8BW/wOwV
mfg3aZXcW1prA3ZpmbZbE2243VyCXO8ahU1J80qZW1a/isdJ7kWDtTCBSweHTRkQw2Lz3Rkdd2Dz
2xJ/ZBQVzzw+I//XD0QA2nlBMHLEvD9bZmMhQLGh+O7ep2G/pd3EUSx5dSIyyx11AjdqyDwfVt20
UXLRFYvRacCoEUazUZIKhEhI2+Mr3jyHdCA5rr2++Pg0tF18ZZHjvT1cWFKF+OEv7QCJc5n0I2FV
M6skgNzFRfxf/NQ+PZARXqbNQA9DaoLJ2mlcYw90xuAvD6S2BpxtICi90NdY6LKR/j/sjwznAldz
x2cwxcIIhPVMqkA1twPYfwFCCxl2jA8TU4TsnSXEIGsb0g18rUlL62Y92t0+Gr6aOO3eSzLf/uI0
vpgslnmFGhXESej4707kPlbx8NIpW6byJd11RhPBZ73NFXksz5EFBU+j/kvews3YvZRRucDk0+BQ
IjJM+GXX4yacbUc3taW6F5tG/QQdEygis/jPTT4Ds4Y9r6Er/lyfPO2m0Z1yH0DuiQRL6061VpP7
K+NOurf2l76ZAgJkMMOXmRQ3PO5R5hpxWRAN/naVyyVOjyJzdMbbFv/UmXmKydquUSYOq6coE7+j
M8jEVr/ByRkaJlcjWGgq/Tq7Wt5iXohpPBoyRemhAdtK5JIB56ak1qAB4D9PhN11tffnxG8M7G8Z
qxikoVtSBaghEnyuvxD39rRazB88GBfNHaOpLiRmY6sb0WU5UOs/S78RnsFD5Cm91o6xIfyR9QcR
MF8rbe4YdzERlUDGl0ayA2G3M4ciZgeilniJoY+TmR2tMsLwlke1oSDmawXAjGT9sPBz0msPqljS
upJnPbERBQ6HYR8IRp3stJE8D5lc+enqrGcXeOxj7KWG8f9jGX1Foa5wUG/QP6jlq/iB8FElPhhU
CGLnGNX4gEemplJFI5lxEtp8bvSi9VEnpg3/c+ib67U9fRW4LCe93KA2fk7p4QoWV2QCOAT3RZZv
rPSDwcWniERqRmhlEzPTmSJwlR9i4fPMTGVjqoOByqXAP66m3bWIK2C71ZfICeyOY2nE5KdooOLQ
L96Imo3XGqrC37qVzDTvjRGGQdrVS2S/6GUjp9nUedFsCV952WlidXlHXxe9Ey0RvIKQ8hpisL1q
6mZMAE8glq/cRkujIXUBtMcLm6mL1QH4ACW5Uin+23QAoxa/4hP4bDX+ZKBYNJGbNXJnWODI0KaI
20wHWvELyp/FaXJPsRtIbhW8VTjI5j+tujZL+YNT5zGV/a3YUHk/xyGLSq7N5lOLe6utpAmq7cNf
ut8EByoKlknO1zKV40c9At6mgF/wru+I1TjELl8U7AndqIuXnhFfCdFU9DbB9glmcyQjIIHKXzxV
o0zC9H5M+Vu1hfbEJZOeks+6zGMq7+eWXk0YyrrngJ2JO0MwqwhhfXG8rv/htjYR1iNALi+pNo35
trrKOZsDaIkFQtQxsrv7Rn/Aj652G5gzuvr2yS9HC3fjl9/ywXOJOmLf8N/177jQ2HtSJTc1Olzn
sXdi2M1jVfKMWwVfljESzoVD4mASzbfIa+s+4I3jZxY1utPDz7q6PdRyY/1vPT0sinPnODl2dcfK
pN4OP1OKEnSIyFSOYR+DeUxf9HKOPA9eZrkgXC7+zVNkWuPR06eUo0FiZPjbBimirBUkme65jkYS
8txZM7DV+R4ZBY2oGe49/Vcr+3xSUzoytCZokoDZkuK1FPIjNE1seG1MY9BgdqfaQLETPzF3fjwq
Jg0YdQsHbl9iWK9h7JZiW5tXDR7BGahdO8rHXaIpVgIFEo4bBn1k7znBDTIPHBH9Rz8ZKbWEfhJu
cpqqIzbl4Asy/MNKIyUsoXR6pPAYoXWyiMaQp8TqH5mGk1eV5I+oeSTGGCELIXOV1KyuVe0CyH2U
3ZtplIbYfdcZcZl0E8EAPbcGztzmsC3ynqsI7f7DcPdYzM4RHLFVSwwEanS90fqltotOoCWN41Z+
jUrkYRhT1Hk5v7eytNSNq7sjVpFCYP1rtnr7Z0TFqXUw+jbmb5GfKwP6PZ/GoGTJmtuMK2HqnNJU
imdpcybftE+qP/+eiDtr5hraLzW7zCuRx/TbhdwKmN9WCix2woKaWjUqWmuPfd1TX7TRMUvJy9/E
QtJK2tfTUb6WNfCJLCd/0ZoUJUBzaXStXA+wZFqVF98u9SoKAwtERwdHadny2RTv+ycN/+W1xeoN
zKSRBUYpLNNhWT1PQI0F5518m1uYUwcGhWed4DHjKS/A5d7wJB99tCD6u92OO6b4WRyCsjgxW2FB
sTwoCw4DY8o3UOcONWbvsVxGSggP/R2+Abs7rHzk1SqkS5KoTbmqN2b0qshB+mZYvpLmTOEtfiWC
ajk2VwF6QILrpMnDJSwAguVa5Ov7AVb99GLtHGxyxSfstrYkf8kZzTIiD0bkdkO34qF7sEJXl2A0
1vfvHw7Suc16beAouPA426BBmEjM2b6ObDFPVzc+cByISGtC6f1PYr81eIwZ3jIW4q00ETXGKYHF
aWtNU/9l71MHokAdn/HuNT0HIapPU5DLnOaRmlos1uGiz04wXYWxls/zkQ8JmFf3fsGJrLE59BUd
qT+BoOYC6tfED6aKp2qerhf0YXY450/gGzSrQlmQkDkSl7yFId1bHMtXMNvYua9ITyIgiEuZAkGv
9D8lB/4trdl7k5Riw0bCbi+leVGDMnR7t39BJQvpv6a55i7wwLPNvoBQxy1je+CtyFUmzVs9oi9E
2CgAV50T9TOolWcj7YVDX+mA/zWTVz+HXh/1T5mLg4QOPwpQy7QjZqpgjlKwR45fobJzoPAF2F41
CKnzdcXJgus2BLYugXBimYNt86d6NuC5L+AYOz6mxVf+TNJeYI/7YrwVVgMKuXYth3YtRvPsBsv4
qlJ0KgeZNEdxr1wDFCsv2WYWtW4vZxCY+mhiHu3OxRuPACFLfiLlF4fa+NKSA62DisInxFptZYS/
izHV4Hw3UloE6WjHalhtPHnipyrfMtQVVtagijEWWw3NWkk+yQFn8uUHVAVwVyjabUdBnmIzsep4
7iqydYmlHsWO0N3hBjPWX0tKQJux4vcYYFB3xXmkgFpyfX94HI+YIHEUyTfVcJ4/J0w/Qy2SjTZI
gqn9G9uHgZjE1heDTIQEw/cMpI2AK5HxACdgoZOlE303WITxY10821YFVRZtw+V+ZynBA4dWl+zN
wYmcQTCAtK19jXromavL0JjfHcQZPRAlOd9Q0RYrH/ww3wp2RgzGtVCvVkELokjufSeGLn2Jre11
loS7u94IYcYC/CTLmrrSF2LahfSOi4/ZUJ43I9fvNQ1rCmojUowRme5091opOm/fgjdg1ESmLdso
q97vB4DJ3LAToNxlQeJz6AAEcXBRU8DGMC5V5gAIRMedbGwC1GOpGbkHXmNY2+uLB641sJBAgBvH
Eu1Mv2UXtYYnu80I1J78An2+dik4uigIS6ewUjtdGptWYCAq6WBUqs/Uon2veAW7taj3U8DQML2L
B7DgPx0955XAdYvZBx5wG0JrDsDoyUSR/KsZivm/UJcxepIWgrvrUAYgf1z7Q28jEeLKgpKxYvCb
YI1kFm7euOjgrP/VUd0GtaCuxx+/AOv1XrzxgLAqJCvMSR1O6BjvxoLXWA9LO6wo9YsyyK7QAzWk
wqtftFBOzBEF0YIlXWqVjMWyTaEb3kjq6dirqXQEIJ4o3SJ+A3TyFkoJmSfsEqtxeCyhqGtWMbJj
L/fflzyoMmKhoDbRj3cHoh6XBGuLtVzDEzhKF0ldE40Z7JDMGRUKG38ajMu/vuF+o5ws5hLWlUAa
60j6aSHlaiPEe1W3NdPdeTnHxJac1Guu61igKBx/OkWxrtqUOhhURZv43FX6DUUOcoHc7ZztYH2C
1HyOEfIycTmgvWFAQmy10j4PAZ8X3kx3IsYn4BqwZtxx4tqByNEz08X8tnn3UQGhw9e3UaTtPBjw
tP/nXmfYQBIQ/CsUXDPdK35qL+dn8wOG6tu95t7ljTq0EBW6ckIKDR5EU+mQjlq+oVk+1cWU+LgZ
RioVsjAagWoL7yYHNfBg7durn2A7znGo4odyIAAQf+xdVuNZEOAAoBUjbdLqN6vDszDKweQVNOKd
rVGp3If0NKPuJ2zBtjSMxB4PCuG46JkJVWHU6js8g+z5L+xiIEcr0r8bhTPW+3ioW2kjeNAIuOWf
Sb2isloci5R1W5SnE0HtIAyFtmkwGdPRSg6Zmszd8vqJbZVbZeD8KrEGuusddEnMtEWNsFMcpMe5
TZNi2yOR2Ath2M8LzXF8PKfpWKJvmbBISy62QdmYh4RGotYlH+U36tUDm6D/PW6XnVexWaKxesdX
xGEfrWGgBlGEl2c8dXW2iFzL9njGcaNOU4Yy6o7LlI03cnjbeJqwl5xvwrK8MoYrdNoLOLjQQsWF
Hi0ay32TFbUkz4TdljRHcA34/HsnPTROnCAQk6cxJdQL4x/7tIb/UkdzjK7j6XSRevWykETQvCxp
97x2ytrDaPSg6bDiUC7/dAxS3pPXlpZgHWIOQ+ULFC2Ms8sKy2Dv4P3Ftn8ekXIIOrN4GeBzaSX1
qJQSIyBiy6hbN92iaBd+Ab/51wtiR695tCueLqF5PGSzRqmXoxDBTeEzxu0R0oCu9jnDiKetin0h
MGI5nK5nbOZWZOh7bRRbZ7AHikKg3dxuut4KLluykcmI8rZMO9YbxRuSat+jI+7GlRncC52NwmZf
5ESVEpX0j+CpqdhiTH2dcYyIfnBvwUvKPRSRcbg2h+agc2BiTa2Q7kIPQkzeGQYOw/u13Qt+c1iQ
AYZ1PkXYMPNVsjsGy7UEguRVp9GBPsl7gn2FQjN/P6U/uICsyHsSjQjf7Opc+xlu3jidhFQhpf/j
2orTag4ebFxpuoXzVQv7ZOvCPU1ee5OlAe6hrzCrvp88yRKdbxCjZL8JHnpYD6y0TX02WO8MrDLY
6wlL9Xq2LHeDdvvWOeaQI5qiJrDi11pb9pYm5nTHr4cgIDmsPnGjk+WP7+tA0KnmbKihwBN5sshZ
fGFxuhzwSjDYeyEnhHFamHbSn9J9NhL+dmgMTM6/6AFn+MahGf8eKY7IZkANGp1TkpmaFYdJZYm4
C+ViUGuAs6ZmYMjNrNoeBSd8mRTjYLGKUWTCGll/mEZorujMrcffPONdHc8AEQFAki9gewEEQR5Y
NWnreZZD5MWsaLKSMjyY4upqMkZWj1vn5rslu4LVUtAl2cfhR8GWTesuPxAQZRYu5A+7prKL+M9z
Vn7EqCHgo4jTz710LTYsTzVBWibhf7W3LEBqyjRPWbsqMov7Jd+zjml0ipACDB2V5TlSqqPcbcyw
meMXuP1RbjW/nGnhhj3BnsVrveambzWpPaHeb9aYlNl1a53xuVgShYzCBl0iMPaoKIcQ23+fpIv+
FbzoHIp99SAXT/p1RBjSBSpMRKghmJ72v1bG11s9fmvfcWeX5qlUKXO1LuFq+ZlTu8dP0pGAc2a3
UdhcqirrpB/rMo95ardX3OZ6rNQeoufqPbZ1to+yTkUgfw1nRxp0cuL9lGunUVjcLr4PA/5Tbywm
sjEKnSpEigcW7fJuhPP0egamh058zdzo9/FLp7jL/oa1LZplT4pqw9wdyESZY9FzVyo17cUcAddk
pGhgLuWeu6L1MGhKe+QVDypUVgBWmWFM+3Ek9SPDSmiGqyDBQoTJdt0XxAfRmx0QJEKMTUa3oPB+
NQPKkqzjRwNbsD1c3gZWQYcbQbU4ey4gCs+JkJuG3NFSq8l8tdEiI+SEbYVChoHaFihiWl7UuatH
o8/d8WbRz3hOpdeRIipAyazc11pFXSTcxkQ896wLN14GvbV6BFtJ0CX2+OcfnG2a4s7NBos0usMR
vCQgg/+cZYzmx0CZWBkeLfGcjinXUolBlDjy5TT2aYQESiS2/4qjM/A4HJ8HrGDv39jqui+n5dwA
DW4NrK5WCoi6cLA/kOYDzdr14LlxBOGtBqrN25Btb5+Is2EYnKPW4hBPhLtmtWHg/Hu/hjy+IUZ7
eJ9TChUuP7KA2L3ECgjL9vw7cL4dq55XSZkbS56nmtaTyLnBpOBWjn4RjaaGjzXiEhidWl3gy0iU
PQ3qvoIEbuPRFUTzjDW0cnBcHDOKIBH1TJ34nkeatQTZ2q5MhB1Hg1eUOzDrnNhekDlnzhbICI35
kMuoEblsfa+XeNR3J3s/b4vCw+itMwUT/ox+GdZzlly6bfy3JLYGnySt/vfFL58Sr4qjra5uYo+j
NjnwDfEgYt6iNEYjUzx205Ea4eO7Ar1/lpwPILU1S2oeohwgC1B9bd1+RSS2dAcI4K53O/491k+h
QIVnMZeAdfOqGgHBRs16aXsjQ5NYx8eM1fuWqvLjVgK9UBw3+/frbORDwp4lgtQGZy19teK/gTC6
IiuU0rSHlsZ7A7emHl9aCEPidl70gXFx4QFblh6/dEtQmb66wS7SSoKicdobJm99/kvMShIooDW4
oAQxWWcSyT+6Fm1YxbfFBc1rcumFbQIfmGvZTiV7cgMUtQUzRAkIFxSjtdLBN0JJWK8qMbCnIvza
skSU73O3TrDuaAlVM1NnQ9+EOE3Ckb4nTZHYyvyUusPq/PRczQQYCGjRhLe/UKnfSr5UA66oAmwW
ifYor6x0y5ZzXMoPNAEuxYYUmcyAGaTRXTT2otxZMUtWOS9Sb/NNW+OAg0hOlIRYNFKVCKmrKVIL
GTMZnf1FXxdKeorjqzXVIxBZugYaDiIZAVYrmvx9E5zCjAQcuYGZRZS1q4ZT7h06BFmlLQV3KZOr
w32pF3l9KLFoW1900c3C8Uh9RhxMe8T67OHAhExO1dnjTDH8gNqCaz63KiBu+hr8sORKdMexQAVN
v490sLpAe58so1cuYdoshxdDlUQiryVXaz+9ZJVByeOWQXUI7QXH6zqt9wNPJ6qHif9GlrBf1JTa
Kyt7sBqZHw34k7c/3E08STRKPNmoo1Q5HdkE8Ho9QORjWk0i7vnNNE1V8KIROgKwbYaRI1N0mSgQ
4XTswL7DxVRJbsFv6C7z14XM+4dGzoP+9aUm57UYa2/VjS4Xg0eO6d2dIfNGdLiW+tZAN2Dx9lvn
XNOo4WGVygI8R2/4c4GPGIhKdiuX8AGvPDnBNlsK2V2mQu1CD799BhSXCmE7cLDGxOy4GDM972wo
XnLj6UtkrimLCqhk0bjb0eAMoBaTw0GR23dZME4h8s5vLZCgq5BCUPDlfBLZInhx92yoEIsW2mia
0w2WCaQaxMKg7hHF7lYcwW4AEy0FGFKggNt6gwzh1Rq3kUjDW6KecF7jJWNA2GQ8QWGCHSGBHjBT
gHtDGc2e+xmluj9hw6QmQ5mu657En3bGugdOCJxfjZjlWuy8iIa75mupi0HAQpraEmX00F5kx59z
yvljrcdcadcLx+3IZ4pW5Q+e1hk/dV5onkQENyovGKD8WMUfR9IT3vERo3KsoDUN/x+cxWpZCb+E
KTZKOV8FLG6f6NkR6Wx8Ta0VYhcNv9Ns6UTgBTxCZPJRaUC/Qse9wz228se8st7iztrPHrQET6v8
b7+AyJ1xEMZtIZZbhiyHp9mPvsUxECcTM6/LS4rWlPwfxkiviHa0621COmU9IKQoh20/Hl5tgc1r
hOnAXNNSAojYQc3dvXsUj1TfZATiL0KK6Rpb5Ybt9CeGi0EbeGLZTDTiKbLkUEdK3zBBDDtnRhj3
wpchof+oYbmhlTQ7eiTSnxvvkn4Os4kanNYdD9SrEJv6Sk4xGpKqDuZklhkgnAhbnb9xFv5aNOOV
OidbDW4p49afP/Vo9n5+btCNPSW2i6bkzEtTMSjB2s+BQtFzzS0tZKFZjWvOtULl705PiVurT/hE
jQV9g81GWnQLEN1Fc06my8GHBnslIroufTck4FXJL2pMpoDiRgwL6LWPmVaJltsIk6FgnpfPBYo/
Vi40FEUFH7Zm5C7yvV0t2U8+LXgwr6YvtSG+jEjT8oSSKLiZZU4FSJo6rBISDQpNf0fgAaWVQt0D
mlRTW+JbXZbuUEKI12MAAW4oH7UoD9t2bQkRnyGNFOoKImzYcrJYyi/szq5fb8r13tt87FVXzW7g
+oa/l0YcvJTMFkfQBUyI9Dm/NNHv9ODevLH/Q2olHLIyONgQ5JhReb8igoOgrwsFTML5CS7EJS2S
OxZ1EMbbXKwqgSsPp03Ws8PyXUfZC4/GhFBxHiNivthYdchHe6NIL1pJQnQnBPuywWTJ6DHuqcIs
vCAzFD93xeLZZbLeEh2xsghetAqpCWPhQZiPSZg2tPp/FeOZw99g6joG6MthDUBBdTDJ5SXoRweV
SSAsLlRNVFziRcKQctqWn++EjzTFuLzUOIh10k5I5JFfAxlmJUMUrZS/rUgTOhlfec/0EVFmlcC0
Hhdh9/Lyo8hf5eXihev/AKP2/+MVgxM7IXyqX+9hfgTLVNVE5rM3KrgaETtY/GH+sESPhiVbU5EF
iVbleAEwHP4qYHfE132p/w652I270YJ0Fznz6nixT9+a+i2K49SjJEf7pvKZO3IvQtK8Pcxun0ez
IoojbafSrKXWKPgT0x26DEr66OFTl//0jIWK2AD5pRdk3pRamOMoEhz24cI2RQ91bMxt8Q3Rvxna
dR8vIkSLD/lLdsEQzbSiJm0YrSpLvXrt3OnGbUiL5LWll2iscSZI4W6khQPBqlUH0o+iefRxFNC8
n996DptlksoYYVnUHO3DIop47fynDZx35idP0nLhWHmLSU0ydCOzcerLz1mIFAJOHrgBxGVP+0eb
taNxTYjjxCz6+SjEao2pwHGgXicfbTcOo59b40BGVkwo3Ym/PWAA8iptGwIEfUFFoFRuq4oEJMt5
hpqQp4SqU7da/sUKpNqMa3mvLMRKgcC0dLXgKrRVK9qgVa8TS7J8U6sEqYXLQYsxuQhEmCtfxSDM
IKHC6xd2qlQZWe4WrtT1zrnTj+Dmq2AF7mAG4ZDAcbd4bf921VokO/xH+qGHHT6TwG8de4KXh1IR
pbRyREnns50+6x7IF1x+ryDfkEsMWOfYC8jgNZJtJH+L0d6JSIvEcmj5nz8Q8f0XcGNN4qTuQ/rf
DYetE1SoyYYPDkBojE3K0z2OcEBFp5+toH6Wlvi3ZvSWE9QqG3rpI0S6HpfraMLTwAc1nXPTIhkw
twKVCR6DlLIYfZgYAinOnl4tLqFP1HhkXi5EiZmmfFbuk/fKTK69WMBet15OslEHtFI6iXjGYTwv
/pYhef89CVkmvhDxjgdgzJJLT271kxrySi/ip7u5OVu2AvM64r7N2RlKJCInriKZGEVKwzNbJ0L/
gg3kZReEOk24Y2PnGTl102fTb5mWW/yipx9BqHyUcT3r8ggBmaA8SCQRcEXCeIrnQXYzSsws8GN8
v95qvA+KKwHvCIMQxywdFim6qIMTtHQQVSq3CkHCS3qU15hJSqCy/ZCFe1GttrLX2NINQRFndWuY
Jni4RlDF9Tfh5CBp8k+cwozzQ8H5LxHnshVYXidIHZWn3ko0Xol1wYmtuyjvWsyMzNpM3s6T+vu9
0BQVVPrg/f24kucN8H6TuVKxNvpU1JNnI5++4L337FsIYY1EhHxDc51bpG3UhH5gmGG84yIuTcBX
PpXwTpcEPe/w3MWgCgQuhMQeNM661Ne6AgWUHDhMS4pqPiQ71E1LPE0qeAUKQkUYRFdabrLKvB4/
RORfTDugy1k0vFt98NRiZzQGFbt68dV4Np4pLhjcL1OITLeJnYjqPoikPyLUPJYch+5+khDHkebG
hmR+s4TpWhwTplJzRnnLU3U6LgIfwYal4ihT8HCMzpqfuj3SUU6IhZSkCUm1zrAUQ/6/5Mb7Os8d
3luVsulRsleU3gyY/qUHAIIGksSqoutBvVDQbQJ740ZBpdeHxOODPxH/SM7VoGxw9gkc5HGaHRdE
AJOD3Z9yxl29/ln01vzntvMu21/UPqU3cDT3ToCTy0TL+HvBHg7Ou3Mjhj6YObpcXdKYUUWANzTv
ohUBkI07ViQ4Ws6BT0QUjHMuWDyqHEH6ZoqaIdM4bjGk6dKUUHRPhC/ZDvRbT+kA675/l1own0L0
w3hve1vfYozbU43ZlQTC5MfRbtktJJHH6rayYiYHOLYXwT9atvnP9xg8HAlsHYkgRc3dr+nHy+zf
9XuRIQYTwZ5zo3+ifuTR0WYiCPCJnoNw/n5ZGNsD7qUZNuFJzq27LqtBiciSDe/rheLnU8j5fmB8
gtfcqC6F0BO68gKfMMrJgHwOLE/Cbs1Honi4kud74eVbt+RL6tpZxg9UM0Nio6F2Fu5G2TPExOzq
FCtFbN5CJ0CQKJRZ0Asg4xpNvlwgarEvC6DOt4B3fXUmD457G9d2zllvg4dTJc7R5gzrTGnW/HDj
y4gUCPDsBZ506HNa4slh3Xcniy3c5Cpxb9dZaoprvfnFBtPoZuL9FMAFqdfH6cCNPfghaSoYoAK5
zEcIR/WJW1Q5xuSQlqcnuWLkovv8uIcToIFnci0gaUeRt2sIR4fOZUCOlCKO2in5zaV0zfJGbFhD
Q5EclHwr8dO4qIot644B5ovNX2+ZR6Y8M2d7T3HTrxBNlIGush1ZC3Scz4/muFPM3hnQT73MDB0p
5093ROHkxakRNnCWWOGeWfwvfbclmLiH9rDtcp6EhVgJCMYnME4v1IrQTrweUpkXGxKSIQm+kJ7W
lDjAajLusktHYq9Nt0MX2yxUC3+QNAGY9eZfNHUEH4Gz5Ja2kj37reLdyOzj6idKDA63/aSm7pnn
HXxnQdL5pFU7W2/snihhzo9EQQ2pchjl2YsXIdyhc8ZNwVboMM6ubA7LiJ3fc98mOOd8E2AiUyQ0
HdERjsa4q4Ulf8lwix1jMSQzsK8Dc08/vuqQePAwmoCZUjBhTL8NotQ/ORU8PhajVWhqCdy9ZHTz
f8ggwjyjN8pXdSBJerTBHWaakA+U8RmNenixZ2hyZog8j0e9XcSmvGg7Cx5NiHFCZmsXjsG0ndhV
PJEEgx6m2EFhyGTkY6YFwfGWa4IzQx1lGqMoV3wLwvPjffq3YjzKrG9Vh1mGL+V5EpL3K8HyHhQp
5e/pYRDcoAbkzla4frD+E50ZCa/D4/ncDhqLOOdWkpvdVCqeel2IXKzWrzxhD1GYEI46hjrXv7lf
hf3Wy6si+oBVNBJ6bi/NhrdP9xGiUl0Z1t4g5jz5WcewaWqVfHXGPS2KdaBGese0K0XIERDar4VW
1/ZvEZHwz2xrqc54gmLTSgvMQYjMxZa0lYEGfIwcq0qCxJQNYVvUTHhlg12HqnfPiNXB7D1Ln1OS
A0F74SmY0SWSLTqIMCqvAE3R9j47F7BlliVC0+waNFoPSEhKpsBZCtmOAcLXLAYFh61H+IeCR/Zg
SQgeLNf58/jXsktntSPzvv2dVJnfIh5Q5ZoBQMwi8FHD+0gq59bepCgWmYrBHFXsIWZhSGYzDaCU
obypqh6TwmwlEbSIeyaTVfU9QT1Zv/1HqJ6w6flhNpljjvUZvJwgTzb3qDPspF3M8VnHqwVtFPL3
efVHMOMnd8nzZBCKM/qI8WSquGZpRZzR6k1jRsnJL14nSKU+mAWBbbtnE+WLjzNi5SgIyHLS6r8s
ngN4VFmcM03H2QWRDk3wXauKP6FccfmNxqkzN5oGAITEIpjh1TCkmmVNr/idDYPrzbvYXp5FHoxp
1cO+15ywVgUWUE12HAidL4gRNRKCwjV9+Ls2PJa/2zW3WYAj7wvLQw972nz+d6ssROBYPQk/fYyS
0uVoqPBgn2VC9eW0G7dNPEwjN2snTHa4S5mGXBANxDBPtFUyugrZs6cVmGRC2ibF9+PQ9l/BpCtM
dyU8OvgDdwDJpV/+KXCTfX7/GGzvKFtnf7Sh5Dvke1RiHrG5UnEKG4BB0+PPsefSojEOSlcHDL3a
sq/ae6QBGPg0kHaBrGXRgGgSPuA471rjTPCqpBDxSgkMxc6rlbOCybMyYxk/ixWqBdyWtaaZLbKN
Ss/EMM7H7T5J2ad4DO2c/H2Rnwk74PcofUCUO+tpBNsBSAFEq9cdPrhlpTko5C76dL6xSLZVyoH4
MVncwyxeEDKxHWwjMvl33Oe27w5D+PC5yKwvcObe9QKxgVB7iwyNFbBlfsOjgkP69A8ReYKV7x1A
QjaxKUOamLpQ4ts4ynTQa/vlcOjuko3MyDbxJBKRfEkQ7GrD4LgIcyytBUCrw6QcW2trOdjf2KJl
t7pA4r0G8OkUEriN4q2q3jHWTWvnp0suVt6Rak9j8VZn2GQJcsp11Oiq6Dqx6ztJD/1kV0h5xYkP
PK4eoWWJ4FUV1/PbuI3DINPqaaT9LlMRUEtW1Cszi1xh5juVpw+y1Yrh+2JXfd/R+1xrHgyZzXLI
ZYtsZhtFOqCTP80pCNDKbVSPdwGEhZ7MCsdf/LWvm15VZ280RDxvriubU+82rNYcGKKSW/CwjBqe
YZxrs3cTqR22Ox5+e9b9wIu1MPgqfP2dBMJXpiBbU6y2yNZyvAvP+JljLcQu0TNl5O8hvV1HNeL8
L+k1Gu9oknWh4/fpsLjk3K513NuBlw4TG3M9RMf5e28I4y1UZuwJJ3sLQ/YKbHCW3rCW0Pn3QhYl
WirBLHRuP1rEP6wb2XuZv0qqWFBUZEpcgJNKA8HvWxCfbguOIc+6+I/drqYJmrVC5OaJpkvaLdi6
ovRCmVWIX7FUj18gWmq6GZZGRbV0H6kDYPLVm+Dkqrke+SVfDcXTu0YL0v/LUUgWeFDe5wcjH9ce
P/zKN4luUAFZHP3h7C/bx1t99uRE32IBgO4dkjrJePtn8YP5UtiJPp0iqxCcAtWfOD+FJwy+uEIe
75IJ01MjmdMCXIAgmnAnz0SpIr8BaE3XrxVjLn0w99DIqJAxSA4/bHSJ3dfT0GWqmX1A0kCx0OWy
A/bY/yKWe8+4akuupXh/fNPly2U6tQ6E70bVVXl9ASnkUSNnkZd/AAmiIgaknF7Wai16xEIWbTr6
Z53yLaRgIMbXhFfFdBmj9xkSKGrtLtf+YJVedDxYRMbHrgRj/4t0tvywnFtQSAWxd/tWgzXTt+mQ
FEvK6b4T4sjEDfDNC2Fx+rpfXtA/uMRFLIJVF/N1MjZucWE5xMA6cH9KHlCh6BjiSgR7y33+dPW/
0ygFlHxOgyytNF4eyZ6Ti7sN2JQISmiVxhsYlqToQIWUL5zIjai++kZ865/bKEO8OvhE2cFYVfWK
uJPl/kEyCTZFEgSRAyGPQVWIn59hMD5Q9laO94ch39zfXcaemB+2AOmSI4ON1+V+/ZEC2FOXJpiK
rSIwCPjq36PZ+7GbjP6IbHkqc4G9UuhCv0uggLp6HyZfMhr7YDqovf6jmbRblxFLiBfJUhQeu7pb
coEflFsNTSabiB7cz100bhoqrhulpgzU5ChHQ4eTXKQ6ovdBCgLu4QF3CELg2z6wL+fyFxxV7CX0
8P4mT7C6FNrQRjnKCRXewBqPq5xme+f5JMf8uujekTDzWoVZTixFf4cOjlRyP3Qe3huxt2lytgfE
JkRN62ApBgroIcfdadbtVtQZkXDxjbtBCluX2pJ3GTFIv+a7Wncnadl7tZHL3YNfq4kzrPmK2cbN
iHEUq7DJPn7VaDtPgXCepXgIKNdZAuTP0vvDX2uyjMDynV48OrYf32dCoyG36dhbuKkysPzdxkdC
SQVOU/KltwQIzFxrgbVBR26Ztrer6bc5jrMggbKHS0V62p7HtjdD4ylTq7tmm+DijNvHmFNK8N/2
VT58dbR0EGmZcgjcqn9Fvu+LdTkXTa5xZ8OcDoPn7ewej7mptwKjnzn0llas89fj5tEDf08FMLYN
V9F+rc28pfGoXpdLoi299tQesovK55jYSYjHmYcdrsbYheG9rnJzJvDkOktfgap+LL6bcCBr56Ua
NNj53+xfwwYaUl6rikOQpyiO7YzorSIlJPcDYtC57yLBOK6y+l2qu38dtGxZ+xHYyMVGCtzCeuDk
NpbFfAsyDqLqKXA15SEQQzxcrkg8LjU/sXapRo7Vw2ZkXn+OsLjzIWA3zkCOGTb4ymPPJvYH8Lr/
0KdOGcEKLuUCQNSrw6jZIDue6higu5FY32b61wZzp1kM6L8YVaNXLC/hPAVdBvhUFi5yY1PqqYsi
IEKxxj9RReT7xl49sk8hpdv/lvycgqQ/EuIUzVvFa+7+n35ZNjfvryjas5LJyBTF0/mSOcBrOFvm
giIv1n0hrBPmrqY5LAxleXbj+a2tgeKm04N0kBpZc5+dcYxNKhjpbb9kYlvY8uOppD1DJPv+P4TE
4x3o/u6Ey9BrvvdYFfuB6+KLrvKyDKdFTISRwnXL97n5+DxzNPC7r9ab+Te9pLcZT+0CG7z9MSU2
Zqkpf2w+35kNXTYLfOyHqrHLjM4EvtRBnTv7GOD6GpSjykYmLJjAyesSP+SwzzWyDHh0SKThlyHH
dybGoeHHFWUQSudIj0ecXexl9miqGGMONZDsvMwF9ggbI9R4ux6O4ZC6xT8l25k+Otgpiw1+wLWA
8WV4UOgSwH6T7JLJhjlVuyymrSfjzs9Z7YubW2PJthQKpNSJ59CBloPcGEVzOQU2WlfMHv3THMrx
Ysqac613uf560fBQZjUKip73eQNpBsXEdRdigdaBnvZbNdXk7RP/Yi3HrrDIN1Y4lBzhei6G+eDR
aQEKn54LYAvQa7ZX1AFoYYbVeepd0zPItAfVGqJbzrkAdNLPQSxsW+/3bYVbtlyeBaUnNmUtqfdj
ITWdww1GRPi/yzeqnpmI+tt79kQmnV6YZj8qwOjefEd5v9L/DAj1RvhfQ6nlC+oPO4jTveNYhcGi
591LTagxInysecUv076JhLy0WZh4EoZFfk0Am2nypor/bMHGqf+UM2PeAgpnDrHIsfozfqnE2nVc
/qQsEQLqm0Fdlkxh1ffQE1smbWx9251TBfN4Jp0uRzGjJzNuIlJfFZwdLBEipCh7vAhEKspQ8QZJ
uKEn6Pibx6kwVJfqzhPP2shs3K2m+9CGSrkPk9wOk1voYGQUSyZ+aMI4tbq4G675RKf+7k4STqj2
zg6BOSBTNfCsNoCIexHo7Rwr3o4OoxRCwkxN9fveNtnMRzKNhhTsw1HXl914lNGdCHEypR+ybTWt
hQnJtaovW5sivTg4df9VQSwNHtRQZ+/NYwk2xZYuMJl95Bx0H+6iNzaoZA9bEGeT21JHzRCcFud/
RyhOU8rDWReidQEAPhny4B27X5V5S57tmgzIU+WdMdZKL3WA4vxtYdSL8nuyTewTx9lbWoIv5/cC
+usZng5jLnEfsc4dDu/Nw4EzWISMOX4Nz1l95t1ioTyi4mPAn2W0VInOAbICMy0TkLHwos/9oDlT
OuvBgeGw7fMsdPVZ1yZMcuvq8noErdYb6FGPtGe5J2X3lUHEcBV1oilvMzE1MJjDXbgGSplcg1ds
Blog9BmPdW7eyZBPxZIOvbsBj+NRWhxu2f+fxM2bYLQHLGa9l5muNB24vnRRWn+gswvYqd1KHfSl
8Hce/LvSPCoeuYvPAuGt9/h92Ev83JzX2EJ8PioHjb9O+RJP0povVgpKTGQOfTKPGMKrP5GICDGm
IrAk5sqiSEFbCJImHhQM8k1Dxp/j3j/jvSOumIsh/+Ufjd2JRBNlXHElOviXAzZQwiv0g+SnLBNo
GpKrANK4gQOYI32t6eEDdZdr4pBATwaqI6DYU8DrrvbrerTV7nssiAOiTHjBoqakZf2pZvmFz9DM
Nb9P71mJmqSULyhxoraviQqX95/CPFl2q3SuGs3KuEwgrx6VGpPH6kZJ1/ui/CRCC16BeSoDiRrj
LsqXk3uAxQmoqaI42sdmAjWuH0MHtBLq6QAkGniEl0/AfN6Xq6Jyd5SBnIP2WXlDSbiUNdKro/YE
LCsBX0lnIW82l7KXEXsGIwChPgl0lv6AXKEgxlrdlP7f3qKJY1X65yNayYQzx+HENQo/px1SK06W
uP6MJBeHVa9jzkxFtSHYZL6IFCCKX8iSD8Rzu9ZgmM2w4cv9vntj7WuU/sEyD9SwpmL1yZKWuKse
GXhO78u/SQyHBwf2j7Ev5PXMSJuetQpQF5E2Q+MJ2hdTQim0khrQjB2Z3UomyV5Yi7Ct0xuTe6Pu
1JCfnIccxMIfJbGoOylLq9jHQkI1At1aJKIpHUH9LhnoPPK1fyxj+jwAU1Bg4N4UIh1ZyKDrisQ9
MYJbm4IWjrooieIB3gMlCHmJmksTCeMs9qA3XDruBpCWpq6+l4ALLA7dJYDJY339N53dqSvaqQb7
AApfAsUGSn/U0YmPd8EgnXM9RqCg8S0uhNaYy7Ic0yi3IF1QJy+RaAM3Sm20B4yodur+0PdqKb1T
o+rsTnFhxLfmw8hC6KEulGQmf9V5YGHdJN6TqgMfgQI6V/H2iH6PrWHHmFkZW7Khpmof++AnFkEI
Ioj/pMmT3KTCgZc+3kxRDMFn5jdHpYBN7zBjAE7ySugLyy3p3HS0nqOiiMC3A4Ti2P/G/JwF8iKL
5tO7/Zlq8mnpVJiSw19jZUbU5Yh75W4UA3V3XRZ+WAcBRVHMUIo3llvPkeHOEGVGizWd08hBAn88
yPAS3y1PneASU4JcPQVe32sKk5ZquTehyyaM8qv8fBRKXVjPyC+8vsyrFOSsXq8Ckzk1wrhOUagr
PfORDTtmVSEZvgXXRaj19VgTXU4HA+iVRACbcqdbOqCR85J+cGhYbNZXmgb2sFS4/L1ZKb2wgQJg
h2cPMkl9oTJEoMfd/O7PVoLur25GRTjuCMgOA0lT4ZTk8AOG1zfdt/S4/xIMUQwjXsmPLYiTgKxF
sD+JshfHXreBkF8l1dalwa6hCwk9syJ4DFDULsP3RqoyQETxARO0GiqkHWbWsytrU1aL0D1b4hEo
KcecqpmKaUChkI0V/jMljXMXfrMELb2NzA+e96vPy1qayJzJWiYmcf+gvqazpGixg1AjNP5lMS41
7jTXm+m0OOdFbf3VP4UD9JtYNPyNiucM6lMqrlA3sp5wRJ+MFsEGv+U59qirwKDcPEBE9Bd1O8k0
wV9wpiX+iAWwRlkgF6ZmHZz6t4xsL3CbFizi7WxuQ2teVn+IcjU64gqqCnlgn9ETPKpciJJnRgaa
6Lm4wYJ26O+dIK76sdAK8kRk6evbiF/i2fA59itygHFNZL6cEasztmXOu8gmSBx02XssiTces0Mr
Totq/zhrp6fvH+pvSUS9qChyLsw/tNFp/rRZGVVG4UaFykEahl6i9j2Pa5qGQMIExJAgEQ+d1EEf
yjluqGtPrvwXMh5K9vxW/fTAytcX4MN87i25B/MLSACPW3wEzuNLl6V+2rRsKL/V5WPK6RFSynnD
++seSeEXAOLdlrp2zWcOFFBDWHrhAjom2Ckl29ZmDRYQ9HHxHNq5s8/Opjufp6ARtJPdHKtZaLiN
o081BqtuUgdeW2zSZxQDWmlBBrv8EE7N6ZOazpW1OZbAXr5T9sIw2aNjm2TNef4/hFoEV5aBA5Dz
DF0EM8Yq7qpCxkmkmIK4N1EXxGwd6MsTx81ln6yp+9emqfDZo/m3tGpljKyB62BeaUe+/mWmyyZL
Q/sxALaqjShMbjeD8N/DOHwiIy16uExd9/P5yuyr2O1/acgMWIzznlpMy9TWgWEO4Hj9MENnX6Ew
TatWJSMfHLD6M6jloLH7wWnVlykp1ooy2mjx10EirqTZaHZFs95ofgKM3sI/i1FZSWf96LyL7aEw
syQqZlYH15Wc7cdahUAcEghAMiJYKnhDw+3G5oXMNOUVUeGWgW80lhhYtih5ktM3lU8rWIt/6L9u
9o5iEQ7YGzoCdgmjjXj+0jnVKl7sZ4afc/8/sjlxaAbYtbHQk+rvhEei2ExBYLSVmJslInlteILs
V1P+V0ck3bs7ZZW4JyJIvpdYGPmilH/40X1FlNnUq8cgMKyNARqFnWIQgN2N4+3+yl4X96z2ACDV
hoUutEr3yzNzwQHQ32RuVHXlFVeIdauVQlLefISSuP8E6F5DYbCNBla0ncg3rP4CFFcSH//jWOad
qAlNgxVP+lG7P9o6/K7WdzWp7Q+MbD68a3IXpvrGYgRbmbTS9sxpRmDW6hELl6souO1A8AB62bg/
RYa+H9b4o+6mcQLRm0lBldPJvSdetSk6aaCxts3GSoWg9RQTHE384fE1Tza+u+ptNt8BXJMHP9Ne
oJ61NqTf+liBHAKnBzpQ5BS2aQJAHK/UBvcD/91AaaKgbYXHPraWhTLfuDZnKDGvkr3wLwk5j83s
3ksTVTRHvFz1X9h99R926oiPwF62pWale/UPcpBM8gLnn5+E88FRM7Y/jExINqU9GHIEdO+5e8/i
5zgf6uZAI4Sgf2c3AS22oAmOY/Ffj/UNn9cSVOVic4FCirk4itqZeXbx6afgehpq5qsMUB9maN1h
VF4TfXtBXruqSmK3j3FWWePuNE64WISukfOADt6sIdRtq5Sy6qVQeWf5robup42sNUb1kfECBaXZ
Ir8z5UOwFPP7XIW4shitmcux9bF/YqhkPPPO6Cp6NfHzEs84CIQTxnMyPOJ8c89QfAzAD7FKpxmp
ZhPqGWGxpwtBewDwiFgTI0eDbKV3sJiYPUwPG3Qe5hhuqNGglXYQKkRSBj3GnK134UbydAUWbIbu
v9+6L0u7X+rxEukUCMv0aiPIo5w2wYI5iYUG5tpewb1kJ/ye6YMEyxvHobu970koODMYtcsP3orT
qR4uSQjMKbRoaa7ZH3e1b2WjzIxA3jJqLkRcWqGVahby3nenmiDxOAxy0CiyRnp+WqSagOoXtROM
J0C/urV9Yz+Siu+L1Q1tfyN8Cc66VsQufyfWvLxRUDkPxOj1lUwMmxBvJD72VJ4cBABCFpSCthKK
4bWxq71w+PsH1hyUpPG6x5HrqDq3+v7Ad4Zx0+STOBy9qBRzKAEv2jy2oGo4DxrTBTG4am1jdm+0
5nQ/Hj97hpKj9Gc1Bg2o1QswzN9KbXAqex8nRX70Q5HwmQ+sY9N0x/rUhKdJgsVBMZ8nEDt5SgL9
HllCPuNP00/bwq4OLkXX0Fm9wRz+l3hTvdrlU/AS3ZaaaLs0146Aqol2dcD2aJxIekhRDZxz6qSm
YDsSYYrvKzpAsdtjggHuPS+7wk54R7OzOykLdTvqcqBm/ErmqHskOSvaVJ7TiHr29UNij6cFgmXU
pbZsBpiob1RH/AQVvvMfIcV7Dv9DAutHYDOjmHf3hzdbWXphikev0C9282xbbvU4yl6lH3rHcp1m
RSVfU9dCWwJ8hluON8oSjxNVOXSeg5wUpgNMgkSg6+Zl3cyE2uMmyVJNtVW1nge0EXEJcrEV+LUa
jAbbwx5A1DnFqgIJx7qVJntSZCgLBCVG0pa0copEC5Dg9Ac3vr5cw1qLdQuwMCsa29QO/FqS59HD
tGbd5CvkzaPjX0sNk+fTjWHrinw9e6SIaMyOWfiz3K6VMaTH6TYmbuAbGM8vdqTyPqLLC8rqdlDi
okHUrH2B4rjfZ3Iz13Bz/fmwT9MsHeZrLhUbNW8F5EkqRV53H/A2zRwi6GIFZJWZVzPIqrzvrZm3
BhKu+O5SUgc4lY7fyaASGClcP5LaHqXCHxKTT23hAFpBrPcbC+dvLpWzoAzPHCz2A8sQBEs34U6r
GtPrfbqOP4WUy1koNtqS+pzeZQG4s21IgLFqfB29QWTRr44/EN6ns12AA8B4mmED1Jtu9YKCqBNF
8B7KVVrATl0nvPGB7mppfhfk2ldSpehXZgRVtj0z+HqiGfB1jPVVXgb3+vMJl9niQX61m+k1Vg7U
RRdXzIUwNPNJqqqHSpZ+WYuqXDlfvVXCdaMpiUM7CMGkCGe055nznW5KEa6kxpNcgCjU34itd7Bi
PaXFQIsJbd0EOatmNvn1+K2gDPZvPf7lFqHH090qKM1IBtyPZk/mW77sLxfbAabf2c9NYAeuc2rL
orNfpG2H+hw8+USD/08IWmk4HnreB3/uQ0Z2UAkFeIT1P2RQs9u+UDQndexrvtEf4GTikkxLsKBf
2llj4hY1ihEm1mm5Lr1NhFqpidnVaknawcxITL3xaNGmRgV1ja0H2VtJ1LI9Q41YywUkWu5zRLB0
KhIDgH0COqFA3ENQaPR4tC/bGNLmg9okGFe2Z3RXfNzDNbum40rUH+1Bsr6xx31SOfYeYf4kA4wD
yTtrUNGZYwNpS51vi5GmMKP/XiCE+0f7BWFxqgZMRh615oYHg2VRCAZQ8ZFinFuu9LgJieQ/f7KY
lUNyx3nxLBzrQXNSFexiDPC3IKTdgu73qvlhHuYjE6wJMqqxTmR41NZjb9QKIkOXu3mTCTbUtFc6
lHF6+4RluVrlwl41sU4/s2sPpWBtlikAZJFZu+9avQCh/SjRPau7jLaziurTrO+SedAOdprPr7aB
bTar5XAZW2YjsEoPXPBlhVPaVYNW9YwFvdN+wRLMia2O35GJmJk8kegd2be0Pk9f04idsqeH6L/P
qpeZf0I3khKGrwTt5XICpFXKBsuEuoUhnbOStBzYR407ekwVE0HcKfltnYytqF3ZKOEn6TLRqZdU
vRx/UnzkjPOd0WyAW+rPjQPx9LuGWvvz/wDnmnObYbmKsVTSTvQu3OjFjiwlF+KRqW4KwXShSfqT
/hAmJMJbWm7faZLqHkyKxFHKOQio0F1CMzoEa/7M97t0zfcNIkByQNn6ed8VWp20QJeNhpkG3C4w
lvDKXfyjzQCk+OgHYq4ncv2V8OVw3gGjEaC1WymR3QyLs8LAyac548waCz1hwv4JX0nNZsB38s45
lmcsPvn2/mYiCP5VtXoj/BnVaDHLVGoORi1o1n+tEVWLvnyyp9cdbgcKVVUJUTYmHF8GTXZKhO5v
3E+tKPmZbjGnxz5CTmxFncV18H3gQQRnt9i7uyefRZBm6YvQ82llrFFVrKuH7iqgTzO37FmRvJsH
A811KlHj5ZcRLrjj86DUXNrzu0Disl6MTybDPsSTg3aKcm7Bco88PrbKk3aPYo0h1DMNPlMGoUZY
rFrnARlQoxuGokz0T3gTR0m7AnFCJsDqZbSeJ6NEmt0/MLRghUnuP/K2WpbDfLnI4E4U2WS9TqOI
69R8eJj2KOn1aWmBrnIR2flLejl/qsItFT+EfG21+iJ80Cti3K9CfKJ5aY6efl3j6IDlGk3sCS4n
h4XHRocn6DkW36RV8GcYj/v9FZ/77b3eBH9fTzhFC9zzx+w9G162/gqxUciFus+0K4a0h3zhgQjn
JI1nfVP+6EU95KvhntjAmURBM3paoOTdOjjE59PtACUE9uU46CJIe/tmWZlVE/9N0KtywWHuVxZI
7gRmFm5MLhzFlnyUSQ6qm+WRs87LpeRLQAwsdkr7/dI/tVl/dZMux1mEWjW/uLrEpPbqkmKr3oez
+/ZLku1sJVnbt10nmgo2nZZVyzTvfXosXTxAoKtBoEB7HT35ug8CeAWurU/SmB+I+Z8xupVWp1IA
fOtPnhlI2klzugct+dX2xb1Kkq9QFbU2zezqt6fj5c4pvAk8ICvDuNV7nVnAURykB1JQT4C3tP1E
RuJUxqEZs7BYkcfmWmTboeYMZhr+G7C9x6/yXNpo6TBpOoURKSreNvAMZ/JxLlzfK0SghCA0Q6wi
lGNSniaDGpD7p4zCpf6mkR9SyYM0c5717nMnpKm4EPBG6w7fACi6rbTj3neZQRmq35991E1LpYwS
QctgvTfc1fcGfF7cAtKsYXDss+8xy+aucEQExZiSFUNnb2UNcPfCh0GzwzSdxsWB+FF9Wy8+yhQM
YNyc6sFTVdUT6n05N0+FQJeY9M8vJrxhxykQZs2jQMeI7VLyONm4mBMYYr7dQbLtJZLYsEYeAVF8
bo+4RXJEtzP2Bsg+gztFQhDDlnyJK7rZFiNozFszj5fX//ArZ7oWEkuvs0vxRisc/H4yJlFgBjon
tZ4NBmSeFdkUBM9ZoRwaHL1mGo3suu72hi3AIiOnTkDNds16Rc24M9qCFSp4881DS+3JkGTM9M7o
2UNTniqufKEHm410lv4HW7D4sRZlL6C3uqB4VByFFK8SM32lVbVz8/22Zmwcx6LAnReMhz219esQ
mbUiBjvKnm33KBV1bSybI3YeHv7mPtxKEiH1+FfrI8C1Ix4/F2GNVst8z1OfrvjseRHdR03mmPbU
YA2Ae8nfMTvEBoDm+X5dlW43iVCDGyjWDCrRyWxwOOTvz2ejIKlprq2SfZea4PEIxw/6I9IpoCcz
6faMoN1FGqf2gLkm4UmMv6flzJhWl0t0al/K6on9o0X0JhwzYcyvy1oHVVSo4gbLtc38fvDC73QM
nFP9nbOt2kkYNxqvPZjL9IoKr7gAvhDdwzLhTP+gK4mtiJtXrtAzpAL5e1Ld/ZGaIW2RAZ+XonKE
L39/vdDfq0ndrDPjUpj02x6WDFOCXcYwQyYsNYPuoM0EUoONbPoePKsuGHkA2iTnzZZqTgHgVCJX
Ohh156tsw2UDML3iW+lk/yflfcR+DBXSMM9sYNJXqPigciVNz94JhC6582zSDxbJ6Rgh0mR3UPjF
ZEYB6SX2bkDiruSj4bXl0MsQecz1+2r86K47AKJ32VBc/ebbrJbdHSAISKpS7WH8ETkAzj2Ka8iM
cex0oj6fBLSZdEFYCMp1LIbFgyW9omuXSQFo1gPWzCjAqroI0pA1LOI8Nb+hyRsE9K7nEYjt4c1r
YWuswolSvmqzds3cz7grX40bCdAVfKxywvcJbT1zGlANEEmpfanwBTyZ2enyTorFeq7Q6ULioyjh
x5nMnw+2btluMJMhR8IKDZz1J6YLQqajf1bRwRDrRb7UCkIEntPVPOBrE7e2dlFtNzcHKl/hPPZR
LUQ22oYaPQrndk4rFeclsiypHxSPeE7yOlolCOP9+bP2BU3Q31PJcQKefSTRIXDw7sRTBnApetPk
AdHQRI/6fB/VJXjNQk5jBpuHoMpq7RCCEnpXAH/Bgqjznsigd4xdbwYjZ8PK84+SaFvsRcVHgmvf
N/P4ul/iq1hkGzSMOZ2g0M+TFYxhwUSkmNr5mnaRryxh8zT5ZOu5icJz/BLfuJPfDzTF+BVh1oXe
yKi8sTyyepVZDOcqGH5f4MOaftQFtRBarRwZ9z3aGZPbp0ArySWHFCUGSaEImzgB8fJUcrS81nkf
DG1cQBsF7niLr+TZEl8bqxrbEgqaPWeOuw89Ub+r/LcMqh6Uubd661JAglKoW613EK5EjqOFjoqh
e0W+u4nRH5FAY3Z79WUKTOOKKJINhMCn63fpxqJU5Wk5HTB8sBec+BGCOEIbEuj/hLVwDR8FusEX
j71Z09o8KWMMQJFhcDC+XLpsp12hA0/tNcGqoOKUz7a5hQYE7fn0BySo8wahDWHmapleO0hlN7sH
/AjKDWFx2Lk29Z7xsbovHuDZkvdJ+Lxh2fLt/ZXGn8T3mmb4rLh+tVNVGvOg4X/TGz/7VHyGoNW/
9NoKn/a1HtLl/9DMWYduBLADqfrRn9ccZii/DGdgFo6f99Ai6ko/9srIN1ta4nc6bTusTAO79R/E
Va+EyVR3efAv3MrDQ/rLAqbRahrPAX1jpx9jiLx7nXPoBsgDcLdGq/GHDFZD0TnBCKIZyM6JEJCX
KrNBHNt7JiIVDC26ICTFzqkhBblGdtx0zPvXqmEHs4uTACigwiVk1mH4IfP+PsGuLuRlTEORwtK5
HJ805JBZvV/VF0CS73JyAbhX4PHLqfoYrg6AwvqscQ6MdptgrooTj2pvbtl6vkKrkUvFGe7GjdvL
wjc72C3TNVuADdWKNNvX8CSVonBu9z5GajXKjgFheEHvAhnUVdSqr/GsuV7lmbIqPKsJjLPLfpJE
lvkx+jWv4W2+1F3HRrmXAJ5EVcnBublebCwqfnYck/79fvwhVefBVhf9txwM/ZSJPDHDaxGU13gL
Vro4Z9zdCXHSgkDkIkZivruZSeXbep1J/rPow+5pocX5sDuqHfduk5XC9fPEUfjNDMeGMBFh5nZb
0Brpo1TqkYp3Ucm2LMsl8XhpBmwZWlUnKiLDPJTmS91aMucajCaUINfElTxIpXIwUsKR5+7BdNav
GZ3nLW6zk8vB3qLoCIZKl5YMyBxwYp4+Emwg8oW8Hnby7/o/dFwhVrOseSngqlMeM6Avpp+73tDg
lhx+KLYgKmdjqKHzwkkxCCiOm2sxmehKLnOI9HLsyjSmNXxSAP8jmhYxbFz6sh99xIyEI+sbvmOV
Aktr6g0xdAyoL6fjRq1FDU+1l64Ons1ZD34Dpx+sj6PsrdiZtbVeDGeyaowZSOB+3hCEdn85DCk1
+L850Jz5RYFmrsQfWSw/zvGmERw43fy8dnT8xSlyC/hPiJ3dVHq9mLMzwHjg1cRz56xgAUW3dpoq
0JfOrLNnID0Dtrkulm1gqq7flPO7M+VOiF5XUs5+rU8mHQsWO/tiLya4zevcZX4CsS7XrQpshVs0
1vLKtM9jbB+Qy2m3otu+TUES0D+BZNG1YfxOGQd55kpl0RgVBhK7C2MGBHZP73+AnvnK/FC2ZlK6
xclsUOfEkEoJi+JWMNeJQTdaTTJpMyGp+ZcT5FCtEF6+inL5h0RA58WSqr2bs6Q3aYxLqLuO+Fye
PFGq6Hn2joAF/XKCFFTjwre/b2MER0ihfrsJVaP8f+NdWUWNnNfhV0VWIT06IODYykPkEFLz4ATZ
rq19ThuID3yGpq6STT8u+7EwGof3iy7qT5Ob+mmJTGtyWBho7wt7vKPjVbKoFKro0OU06H7X1DDm
/4dJvhgEUT4op4DmMgEBW8eGbobnlOU+dajv7dUE0tjQAmSPmzRnBzEMMSCEiqC8l0IX5JHQJwar
EAMEx4kYA/t6p5sFqjwb6sfkLjL2YRLY+QWmDVE/Xfd5vzN2x4T51w3HiQumj80n+AUnd6OLvIyC
eH9v9tokFRPuN76gWLSU5rT2Dw8WN3h+bViU82aWGqW6ft2or2vS8eUN0sfNiNEJ6mL0ZapAXpo7
PTxOJgWW2keKdPRe6HEIdthTyq3L/wp+riPqxbOYS1tNAHRU03Kl5qhZgowk7BxnEAeuQhu+kZv2
hgDSfsaJjl2Vde9+sMgyjlpmhp+t0ZZcVNKk/5sDrvPJXuy3/LU2WMjwFKDqz7X2ELKQl1gx/tz6
npDokuVgyxXt8y4s9ZhIr7Q2GI1KyhqHI9TRnOKsydSNzkIqoKU5i3rJ3LtRIWL79n/lb2WwKofp
wjm1fq1AoltjSHfaOpK8Dfrp9DAWjAPVh1GW5kj78FVtZc/UKer25ggiH326TKNXcJGzNKnDDtcg
QzZ5TjhNTcU8gQ/huKI77LjAK1b70/oaffRobp5nlTtJFN1U5fqy9wTtlMsvsLrDU8boloLcvEhk
cH90AG7YKz/AhZvCL1V+sRERuqFdqthhJIrvyZOp3Qf1Pe1qsNMOlAmg2uvYecd3xOUbRR2QLLdG
TEdJOljAqo+hdTRHfmoWUXk80JcUG9BRpkcAeoSVW4ZBbSx+QGyWYI6pXg5gYD0ivSkfPRltKXcx
PDeyjKSz/wBrsQs2r/Pj6NytJNYbavsZFkTZinztxXnvr77idRQp28KY9WrkGWHY4/cGiKA2Y1yY
Q90p74GkybavWXWQcyDdb3dkjK/7AF519pH7dyp4cM1/9Ibx9s0qUvZbOJb8YYwSa/KLMxupy3pq
fCrx62gOteUvGW/kKHkWbvtcDF6xyClpL5xDxeYBWPS9rZJ2qq6OzhGEqWqnMdiLWbkarnVLTqNC
1lsKHk58pG4UrED25BKE41phBNxDA+h0XXi5Se8sMLLLyD8QPCsYgabc4V87nN5oY2uKOHVmcOnn
jKIDEDovN+gM4gqbiDjQiZEYElWcW9vWd/82mR1mk5agACc9xeeU5JNRIw61ycGFkklgZfb1Tga1
tEhHDP3Du/kSMNOOto3IDgFFT/rWGSaF5Vd9IwYSejDk17ZInT/wB8JreqZYeokERAaLcmINgyLf
0X2i5KuWFCbjzscmFeRLVYpMtgtnGAm3bZy+6/0VwSRmtoF1eHfvBKvf05mU5JI28rPqkJcv5YNd
im1Y2Bbz/IybqxsboAYnbDu+Uz53Gb9ZBADxicYOoTAPLRvxH2bdkIkivvMDhG2687jWoLcH2JQS
a2HCSBtW5d/7hYNAjH9/Ype2IKR5Jp8lKvz1WbXhCPHiwZ3joVatVjTkn9rTL2i3PSgcFxLSw3Oh
H6E4r5H4O65riMuYbINeIhOFs4ruA9zWXYn0lijQ1U+S1Wu/zkPlAJelAAr1KXFUAI6tfLAKa4Sj
vhcXXccBI2OQcxujUtnhwmrKFs/ppPIKYQWx5R22Kqx0qrOFqFB0MW0vZ6tQnxVlu3hXUPBOZQnx
N7GtVW7tKMH5hFdaeKKWf1NSpK0PriUZV5em13rtUP0RwXSzvj1Nwd0kVOjUWSxp3/9pV65pyKhx
m9WnJZ0UgP2jd9af0g9tIE5mUtVeJnS8yNm1huCjr7+r7CZk+iDG5Exx3ZZZV/KNqj126ASeuCfe
TL9sn2Wc0CGeASvNMhE4YI+B/hrcdfhqyrK6IrZRDwgdRsUbFzu76Xe/Fka+2f1/pyEhur7kHBnz
pDH7gCyv0LmWx4TvRyQfiHH0HJhEjW1o0tf1XQPAqg3zJgwcFW5ihreQZBIgCpN4k68+QM6oGIOr
HgLRSSQSGpWJSdCNtMFX9k9qQv0kAaQr3blPcE9l8Oo9t4GCuvLss5zZkRtphiw8xOX+Ios3pvpc
7pn4we5cYcZM4yQa7a3gVV83kgphykKzrrXjG+BzUDV2x5TbmLQrtJ7uS9OOE1iJfPO9CtP8ql4X
A1pS0JiEnmyklXx3HZy1RKxXDTFh8NQaNsRD8AJBA9vVmN7+O+/T3ooyvAbPgScwUgyE8nVNT0m1
2RpxkFXKLHib37Fkmcn3greXFHpftYqYyHEeybvfMFm+OWzvvUJxlGJkRhTxDLsobMFuTqcjQca5
0m97I9zY/tmDVzLsFB0hQ81TRsz8SbBlf2heb+0EiqvhiIySuanDiD32oEGZiHQxgOInOU/iKDS8
07Xl95L1z9Z0sk4wm3jMjQY//DE4d9NUODTyQFSGK/UPlB6o9F4MUsLZvmYA8OKDOBexgWLr/Y7j
Ygm4804mZ7chCkfn4ja66vwkhkmnVYeQj2dikXbUW5m12vshpShSFPZEama+ak17hB0paffS0abU
YUihMEknO1Hd/TiidtjTEtQBl0NZdr1kIh8uuelJkZCktKF9kTYiprMZ1/eFGzwXHCHWOiT9HJgU
Ld5jqmB9N3jZFmeUoqt+Me/C3c9WcDU7EdN7+h7Nz/l6+pEtPi+HCOtZI2Z23X8xNW4qZh+8V8v9
kWEgGjJByrIrYQTnTkvuJv32UT5qu8PpNLdIRaEMV2VJDALMNJHTcY2xUf0N+TJVQhs7V4oeITsx
MecweOd54ejYTad8tpuZIYWVfD3XGIftmbGvJI1LYi2MH9wNXaMMpFLI/6FxbqcqO4RaZ5shlnEb
hNRHhC8BlJO+8yvm26PrtPBm0ZtRoWfg76sCOdZp6J0zRyU/yt19r/vqAFbxTWfyfh4p77Dzu6BE
pgdy2Wqi3/nedFYB3sqtClLDEPwpXmzDDb2SdeXRRwHSwa8Sr/HjLZ/y6I/FuJXjAqHc2Yk53Nt+
WeUheugdbqzsXY/BkDuoB7B7efsZBd//nvXucNS96lE2r+o3Xh/BYDsEImKvEGU89F4DlzLNaQWK
TDuj3//NPwvOqP3OPLw1dI9pJ3qdEQR8pQ1GJG1M9CKZiaoBtvWI8LUtLZOqF73bDTbqfXG5PLoz
I8/XcCgWzS0j5I2r67dQ5i4M2d5jejfFgFykGFBba8desxLrOPo0z21uaWPFTgJcmxIojUsSqI6L
dlubYrQGOKw9zwMD7RGZT508Vh2r2JKFglrePr6Y6199B/cqIPjXlghJd7w4ezp5bXA7HeDFuGIl
2S4sQ1CGmL1VKvKSPjvvmPEfu9pGZX+hgWQBTNxNme7xTRtYFY0sd5AVAsWmHvbzb18hxbqnNxZo
1kyVrN5msnw5Tyi/nngmkjxTOFQqnAlNKhnoVf0GNSKuuGcX9xFUY/+TozOjYrI8RoZIM65oKuF9
vJHCGFVMLWGDSIp8WInrBgkUht6pniRXP3LNHYs3wNPo9YypUXGSpHcFJLZw8Swc5dXKC6Lz84pe
MgsBrZ6kA/Ul0qFJZQyCAN9xfms3meETdyKvQhVIcUZWPNm21XyAgniKaFVLX9563o5yEAOtNdp3
OcxT7d3bMrWSv6ekackRdtAcvrO5TQ0OqX9F0AqsZs1N/z/ZPrCbShA+gB7FLiUE4Miy1e+IbAJ/
eyHk36YdrrJJd1l12Hv8ehrCIFsOG5mDQi6v24j7AgYItdiSkJRbM6OjPbkQP7d5UGhiCNsSLTqi
z0gu9Qz0/ptfd4uIA87z41qT7PoWXT4mdUJrZ/fNeWF0hXtleIYknnIVEjnR77QWds2cyQJoVgIq
Now2/w6j1LXLe0yKi8Sk1jU1hsUuPNedsIgebXxtVTsj+iiW5AynXf9jW+Yjw7NpPSvL1sIGja5L
ZiNRssoXSB7XrzOdpNclbf4mZQAEv7A/Gy4y8C2xmx3tjScw2g4pAKVZykjk7bClnN3CzIn+3Tj2
r9DzRYgLIs20GdZUZJaB1nqJpC8QWcwmFkK4QNEh5M35+xQCLXHuv/00X96S0UP9dKDDObLqNBsX
iU2yPCDHeHlf5S7/kQO2rG8rLlRyc7+6n9T4Yi2gnLApPw2SKyuWQCsBGQp1ar/uLhNZ7QsxgEJw
Av6ir/ZPkOJYNBSiFPzVMEhCGp7cGHrfzXqc1FzcbPtm0sSC4fZGdVK/wydEGpy/RTgRwc33buCe
NzZe11tkC0HstIrGS1fRX7y7tiiwx2vAe6dfDuisUnysyRMogrO6BubFc5nvSC5/eb0UNGyERpDD
QSLx1+rL1M7V15iWmRYYIHiVvo5KG1p40/CXA1LZpUdVUJ5xb+dyN9BfMBGHGTrMItY/3vaP7mYr
g/g7TfhYIN3HwtNlpFbdXDgQs8GDM8gygRBZU3+v1AWuXIG4eR1XJ5HaguETwWdQQDKv03y9I6N7
AAS38GyG6ZJdwaeioOBpkRytY/uPl0n7CUvqao6V96iqdw4i6Mh8mMg9rF0KHDztuWcO4n2zUpfg
DnKFVeNbs7LuY99LxeHmdoJQ5l9pp5pCT6Pk+bWBOvgJds6FPBEFHEYH+xi6exeVB5BSa2cIc3uG
s59fCdMKrnJTjb89kh7lsoC7MOCXQqD7MaairCRA0+Xj+YzqC0U4ZN9Hyj/KqkQSpOaMPeGQc4+e
hDuebg0ydGHQVd/QgUnFaXELudQQF9k6VVw4q6sDFA9kUm53UnmxrsdvKWPO+HCbUl2RZG4C50f5
RNUFOjT7irwgFdqXROPHXU5kUU6YprLqUafePI3mUpT9BD30iw13q1B5R2jS9ABjfr+u70mjm3pQ
+4US+RIXVwrOSgODR5/sTWye4bl08UcZ3Gc0Mf3QlM3pvnJiwSxsJBXXB77taImTYEjqvbqbZqIB
ZXL4I8/NOH9a1u3Cn4lyrPxiwkBS+R6mOVKtahos6K8LPL/lSK1Efbd8lSEytuD7rDEzqKdjrrVr
BooCoiUMa8FawxMnacNcXTyEajQN8vRGGsIddb/6iDg3dYmtPZJ1dtagKKA7aMW7V6mYFj4btV3+
Gd9G4zmNczmeOVjpo5cQvgl+Nv2ggBkfuWR1DHVW07D/xGEJhs10Rxx8rCETXK7Jo5u0WmRX8Tur
K0wRlnM0os1jaQ/BFa2NaHsT8cxOuoCIDov63uy8Koifl92jUtZrQpagLZyQrZrRfqFqlvFPRICN
MTk+iyRAAWDjNIAOF5XC88eCQijjEMLBA/RNswpWwDEy2M/81KvAM0QNtuspqqexkvfS9e6c4Sok
IArVqNWGef9Pg/RLq+ujU2baSRIaE4fXctOt2//sS2AY0UPXL+cj88TyM3WHxXP/AW/vkC5rysHK
VwOBD7KCT72Hj+wqmJwZnQMSgA7nm1zKs4y0Wwfh+JH1LRhLmNZ1UA/ebFo28MYILCQwuzYrjusa
0TNLYFo1xOQle2CaIildC1SKpcOalkYsg8SBEEVOReAetLM+TusdnH7gggf6RalY6oI1LEVoIkXL
BCSOpKN7UJJs9/21cjsb78o2l6+ccmARHkwyT7hoQeXo3RJv03GFFv82Kgl+4oQALpdfpAgK20qk
70nztx9kpkETAwbZin1Z0yP2HmT9vZ9YZEypCgLc26CZTCBu0pKx+EabNlQ1LEg6uMb74KnPKHYu
ai70SEjIMOGy0VNYLPilUEemIxUPfPCS9oXLNPUAuXkaubfshUU4ycN4rqlqYP0GmVD/G7ch7gyL
KZd5K8mxGiPORn3ua5wcr3hxXZ++TAEk61Zpreyo/7g+R6fN7iSJW51iTv8IJXfXe+ngDg9AiYQ6
HsVfia5cJT35UlM1nh70auyElmIC+j38Y4PA7cTyOiufwphlamBWvinR5IM8R1lYw92EK5h8NWeu
ydlzAEzDeEkTWLsYgIAXuCtNAiOxVVIW0i8yxxvAibrDqIaskHbj9BdMjmrciUuLaAxYU1zwlENp
I+3CIZ45D0V99g4FN2HpkMohqAJVi+3vDF231Wao0ywT6mga0aZfVgpM7BP1qgSX+C/6QLk7FXt+
sutSGjsO5KoFqGNrKYzDYZ3Ur0bpiKOmQ8YcbOUx6daIKbc5mNKL1aoryR55qGVnWrg5wRK5u9dd
KTeRvLS9/XHdCqJQpf2q/XYfnQ0n/mILoaqgO1wOZZLXANPzZBpdnY9lGnLTuAaUBOsiRGQeOeoP
9vxRRIcHsVJwpm/+WaG+XjKmiUkIMuJY9qE0FPCf0fZLPyk5GFT3xEFOmXpvOUGcM2cNC8knilf7
CVfGaHhml4dtS6enE2x6/JOvhneBpW4RHJA/KYZDU9hbwaKQ1dINU8C1Zq9+ZG12OYQcDXimWRRt
/S70uxNSOizrEYoB7C9zbghnDWg1JHcw0lB6N3swDGPAB1lhlZq4+hqfING7xF6yiYhcpLB/snDA
dwQR73t2sUrG8/EBWxjd+7RpgyYkwTrhFeuc/zeaTGaqYumSCohldK/+ZZukBEMbxoIZMnoX3FmG
rG3B1Drc43U5LTKDVPhgs2XOSJ/UI4AOU2Y+Evi9NID9QDW4V+xh37HWx8mkm3ngsj9bimNBsx0N
5FPPLSGL7Kj82q6nujrEjoiTwXRmhE1G9pZ6+IZNWWkmeXkZXn846jm4pwUvQtgXA/+N2VVMVGNa
T0k9X0T5r3yFzaR6/dLDNlT/+EmqHH8fclzbWhvxmGcy3TmVcAubh8Okk7K0Otw6kGVpqr9PNNYc
iqvHEBOy0MXYpiChCMVcx1T40ACLQfWo0nvbUvtaOPzqdHWeioiWQ6kM2S+bFkz4O2VyP5ZNatH8
fFKDKT0rT27EKaSo71B3SYmktRYv1fWnGYzc/OewQkE57nc7y2G3egDwzezTCAF/SHv2pV/GQykF
j9exeT6b0IJMoEve+rVvTBtejsdg/oTGADojZsH7mV/heQtZMhrlwOEMEAdqwnYzCz8EpLOhExO3
s9/pO2bZbLr1KfUTBInweQN+kJog9JNGG/1c22SvvPuyUD6nQhUIk6EFt0lqY1YtqbgRFe8y5nE0
fEqqdSiHGOwEndiWJrAkiZHYAGEMvoWGOVcGKprCdR8K6xO5k2B5f4bRlF+sC4edxPDiyKGVmTnP
iUClohRmbDgNTmGixOMVx0dL4QkPSuaL/dpWl2wAt9kMXPdlKgSOReZwg/XGgISm95YgQElpkQG1
IFnwBiq+7BiUekGGc3SXlW4/3cHSJTotSdblCsspU9nkjkYnCsnslgvS+D0BsgqIMbQEP1ekbpZZ
XM9ieZVIfl52+DBOisa+v4TweNociVUPC91fN43yv5/GagiSN8m2N4KNc0NkL4RRVmEDmz1Ksnp5
9Xx/zl+ft30gXIAivbFkJPlmh23c1j38X4AfB0pKp02NZbisbObs1mVIy+z8SZKMX2F4j9ATKLCl
jCZqgJ4/6PvuOkvq0hfYgdnRKDBZRfkvnZWvwtqGC+k8J7FNdH+9Pq7fGPb2hBdz6mosjMA+zoCo
PI4uk8sViup3/TI/uXUjI8AemK1K5NvrQyCttPeVus4YM5M9qdvAShvADUhtI/t3dyKMN65VVGyp
XJlDOaGIRwP0205IC4aRvn5lAEKKl4RFdMuWtmBqXMzMFVlJ016X2mlVnrupxR4XBySpQRSoEJth
a0k9fRVC5nA/XyIWAur9PFm0zt2ylkB44J0/sLDwaZqxkP2ygAihki0NtSX96KSxhsKuUzYZnnMt
kgMgazJqAl55luB2q5EswDBy7dqW2g+nOkZnFVD8Z2INEtOK2dUsGeQHE3x8SyvOpxn9pm1Uqsj0
ruVuQGYeSaTV/g7b5/qzX8Vd/uz7JgF1Jerwm746AItAikmyOPGhc+GCI1q9YRkSvteF99xO9Eyw
Pdn0YccNVgMNVxGGZyGY8Q3gOUMz4nvlrXKsmicb0tpaMj/r70qHrJuvqZ+pH9z3wGBNAGG+G3FT
OrjFJiYr3h7BPrTU93MD3gF3GHUAR2O2q5eamMPZlGBqvv7OpaZXCvM501Pp43Hb9R/1dYvD5O8I
ACe+6RDtO7mIDVzMDos5Y/uvevYNuWcvH70R7s8zuFHefW1x0BYUp6CqXPY0IzTN9JYu/wf/V0NL
do4LEkMalrRYdWg1E8CYcjB6K4Q0uCObk7/KyShSC0TwRulG+GtNWmtSxIIkqwqzWZGN5sWiUv9a
9PMXPbLxoN+ontXBh2InR9ttf6mZ6I2Cptgi/JWm3sfiI0cG4DFeDbD3LtGU/5bsZmotFiJ9cIQE
uz1lYebas21rr9bxx8F1yCZYQW9rpRoknRAHz9ew8d6efu7ha/iP3C9FljAAmh4zFZddl/GOfP/Y
ep2E9ZGeHKA+ThaUpq5V/MJPD07g8qdfOS+qLkkynlT3XNiErdn1QeXk+WlLjFiQVWeTK2tRPQXX
dAwyXpXbRwsqhVz+o48gsEkaDJ0BBqJsbKBozTmRWAIbGLVk3YSk9YqOAOHdbrZKDU5jHcgPakdj
xpjTPHFx0WhG5Tc3ZDclNBZt5GvSfBT7U9QsbIy1VrElKzZbkP2+d16E2ccuw9KabARNUWZxkwcl
do2hYcDSqPOoODKvI+CGpNcyXAiFTV59mQxoQVnsBGrGKO1ViLG72USNi3gbM2ILXHKl4yfES7eF
EnHDlwyN9AOyyPG7B9Wll0Mm1qQWWkE/tVhWrQDFnv+DRGzpgcTKh9xbAd9bXcEEK3KEMWSanFoV
xyzVBhwITprwnDYBknJfAcRaBAHGgx450vyodRXREpRN/GM1i69jgfOg3ESK7NFP7nCX2mW5aTDg
bHwezURq1cdgPhUosYcgFI8cL13+dVYFYoPZ4Fcm7Ct027vRyG5gKsz64CK/hoo2RCM4iBFsNJ3a
MsAztRhdpaso8SbRFE40fCMiO/VUiL4HTTXNSVHD3Dgx5v1jDjBfbvea8X0d9tZs/fLa+RqrkYCn
dFQxQRzeelatjM6artGt12jB0Juyj4DgFuPgzM2HqhDrrIKBFfZwsyaRUgLiA4LBk4TRYT7v6rQE
ScXvltdH2b14yW8B1K9A1uPXEm/lKqDLsCOuXWMmtz4yL/pzGdr3RuwtLJGBEj7+y/BGy0ERGsdU
/nRVbnFDHbenGj1QirzllNS/lyIyKoj+De/OqPHsDlu8wgJEzPiWF/4VWjgxw45JvM6+dxB+cG/3
GO/DO+2uuMGtraITI41XvsbH1sECKzmcDUX9vfHAWIa2pw1maZwK2d7FkA7sE/lKxzWB7GlSaZd3
sS64p8tB6eM0wx26Q0mqEr8TckIUCb8Jll0lt3CAXukVpZP6kxkg0G7re8AGfT5OJ324oAWFwxRr
tmS5LA7zHuIPsRjW/NW6spPZ0kg+Qgt0T1lGk5hd9IRCLVwRhEmMRnAfXiALc54wwVuMbOnqq5+F
KOM3YErbqJ9UCbiANSs3Ljn51xvSLLRdY9BJBrnoMGHOT5ejlCAWc+xGxyKDO6cAWjKH19ljnWcO
eaSCGU7AJczL9uBQPry/ZuZ4xrxArOpwdhR6OIDp/THepA4Bf9dajS/rL8plomJWgFWeXFEyx4mx
0id0LKA/g+ThWhsUH5266jfO/pqfHHWUBiJyuXb0hQObHPoea7l2O3hKq3gQYTfqQyxCK+n2MVFm
K4UMASpjLGKsdV6qe/G1Be9H6A1XqTnRIacQZBNEtV8ttnt3ZuIdsrU6u1RrbmYwLOX1DeZhBuHL
vrvSZHZ/+W6laJDqHbxM/62teUM8EIEi1/MVEmFtRBSaD+QxE8wFEH8WyIANIvYTWyHIJVWePVkY
Bpx2/8waLMVEYRwW77pQRYgokZLZbWdHuts8AgWo935kJ/BknI9/VHZJmM2Rlcy9IHo6SzVeMJ49
p4/8ASzzVQJc71+8POFRzOEeid1pasaZR389wwfR46FpzGmKXfgQwJGJu9D064C6ihwKzKYqC/w8
G6hbt5OTQHX0cRT3MQ9UWb6kgjkQA8SEgNUC2BvophRxvivziXUn4h27aQ8gfbuUvOTtz8lEdy4o
QqQ04CZVk7uOa4y7+spyfg+OKYHk0O6UtJ4mvEuhJTxdFVrazv1po1HG0bCIgET0JgCcGkWy1yn6
iWCxzflSo2ANDYWDVk40KgEaW7RTVKDJfcNr1+hRahwVmxw+xLfqkydiFv5aUNAO9oyS9J1p/gUP
M9EFsU2n55XK6zllItYIu+jUAgeEMGt2pnHDaRF6GeZpZJK4IviSe1GWKT949m8O4KxeqyGUXiqx
u867KuW/zU21JtM7KYDTczorNNwXz7kUFbtN0KGf7e7A4BbojPhOQyliqNdGLjFxoFcOQTrsdsY+
CoKKsI/yI5Jhhx97YfxkDXpWx7IaZjpm0fAyolHtebX8pj5b1L7I2kcAI/fFddPUBxEiaKFXz6aM
Ml69UmMr+2PfABZvEvk5CeAfESyGQylkLiCGhTcmgBtBT4io6bqV5gi5P1BkmEwB2YkKXV2Q1hHE
XkpJjz5ta1rW+fn8D71bhc9suxJVWagLnPZjHnbNDslyDztaHm+OOl9cu8sIJHQPEzsNAPltKkkZ
3aYHoKN6o/i0a5BrudUi8LS/yKlXSF7NhK4WbDaoai8+HQzwKZ+WfvIZsKmBhKIhYR6vOAJzM9K1
QAkolr4bJc17GC9SNTCKAvCckGcIUDQiT5i7/XsEQLqs/hAKYMKsWYR6R6EOe8N9jdIFMEn/V9Pm
7j0/0VaaTwlKd6GEKYRWOXzMbj56iL6PTp5Z8NPhMzr9ZGsJ6PBMOpNzIf6b43VK7rK9oG+z2MnO
hOzVqhuHZw9ZVoM2Ez3Xkn3p8DE+cl/vNzRWcIfgi10GXVdfO8VY4FV1whpL/HSlHxGDJSA53AAo
mG4fb96TH4DO1TirpJQcHolBMlPh1wFZBDpdXFpdmf4VOu668SpT2hQd9Xmy1gYDcNfcDEMniqQ0
VFubwrB+wIYR1CGIvbu8biHvYJ9lq9WId5zU8pZfxBEtlK+pNMvLpVPkzAWPysa4u+kuvFxuXcU9
JrVDtE22tRpTu29eR4e+KQxuhuChLDiUg4jQ0BLO1jUHTv3DGumfCvt4/dGGwLBmAu1jVaRwksXZ
lQppXPeQyxadhanMfvRIao7x3V2BU4Dflv8LjnkRwnr88beOtMHirYRIq6GNWdvwtPIDqXbqm7lr
x9VhM1WOpsQ2IPOBNVx64TwcnYZlikR7D7PbXqBLTd6wxNU9VFbIFZkdNOpRkMp3uUkrAjvQA2w9
an04Xmisj3C9iYlRwPdouBOWXprxDAro7o4XshAJOTUje8CCQaBlcBXZ4mrfM2HzQ15qDS8YJURQ
tPZ8FqqkojO/KSs8hwLVXEU7UZF+LBwccj+jgYwKaVUTrLLpO9b7PRLKZV2lsClzvMw3NQOZRWpO
nU7TfBoIbAid6c0qIXppCwGWqYZAozt/wOZ0MXye6X07zrEqKDmWUxogNy/e22gYe43JwA2l474e
3sUnQoBiITgyfBbB5PCR5pOIHgUbdCKnA+6iWi7tqbWff8geol6y1n9QNwX2SzPMX1f9Vr1jtA37
w6TigEZfbv+SYo+GVtorYZDzyDLPbQleWIT4XVx07rAYdRNPEcUbI7LMuZVmAsdVishPcKoXKcBl
ds/zZC+hTFecYMqpRn556BQR4n21fNuHya41ug94+2ovY0BrgJAX0xm0uOCIUfvgqYoPYe1MhwTj
Gfj1dqPKlOT/lIMBCmt279k9geEoBU2QnFUAVHNKzXpDPHmpk2MmmNKLbNwU/PkIDC6xWur30w5a
WgVu0G5oDC8abb0F1y1w4TFzrhEKhBbEE1r88eLliF9VaVTpz2yR7R1UtNkJjGjd8mk8LbrzNgKa
hsbNkOpil6Md6DPqKAVxm3NX9YioV9mRiwLdhydAYRXfsSfXlxiyRmjSio5NiV0rPsfDcWNyqs0+
k2MBiYMakdX+E0mqfW3JuhreDicCGTcQ6JM1EJbCDxpeaAnD0nscHizxkTN9JxgcFKRYn55Xsb3K
2oCGYRcLz88KOmqQiaNxCqH7OgFElBwtdYsB00szxnSfIXZErCm336PQEXRFb9hqc08kCw/6tYux
boEZ3dTHEgEQ798hSQQN+Z7KbZi2otTqBMvBoX6A/hLOnpAzvsMsC0ZQjtY3BeEtVL7VciFKJIno
izEv597QRoLNsyxZxxGEhRhWQBxUU5suHAXEQIM5ilFbPvAbwi3i7C30dJvyio9BdDsjfA87iqQR
HvbfnMVT4qTElzxqk780yEQfjDfU1hX5moYkOIuqO9LFgldhonvbdwkuS9Ngg4UtWDPzSO0dipnZ
GT1Ca6+8nbVWqq7lFaUeq3PWKmjwBoGVdedlenO6rScvHdL/f8GffI0+QfbY4jUON63dGarc+dmm
QWTAVn98s72M0seMYXchrUfMkmLWGSNSPP6Djnu5T4OWs8oSCKZWk+yNnhzUEAQh8QY9FqcO+lmf
+PySh1/9rg7lgOPH8YTVQZVB25CE/nVxzl5aLXmotR1s59VfA2dBUMQyYoTMJtKPgYJWvzYtugY/
H5tGy/SluUyA/5kXoiP1yYXimtDjvnk4+iR9iylwvgfZ7mrcipgmJ/dDT6gi9zA/oEna6WV9G11f
p4AeV0wMCoped53Y5Jkyzv10HqGT5KKI+hgS8TO+8eRLpi0KnfUxM2Oa03ckbYpQtlTnUkeZYxjf
AyWknkWtvaWxW1KAgHyC6uOagLgy3WUzhzccisunO2W2kHQE8DQfzgYDKx2v0Ue3lqF+SCV+Sml6
Ej/kx1FQ+RhqEWlcqa1F+c7ZubikVL2iQvVr9xh5iUkmy3gDdleA9+im4uRz+tUFI5J6QsPO+hzo
OSLMEQJoLQaW1wpZ+Zp072XNo5sh0TWsXzr5QtTtZW2gPn+/0xD0heuy/n9hGYcUbM0+KV5KuTku
PVgqvaP+WBvRZRWeOgh8tsjOjvu7hEQ1pzSJMV8wkOxIJX7S03BZhWv5WduOm2AommJc2Bx/6L0P
0+HUPGRScer0SVfXcP84ak6eVKEwpW8mcEaA+hMR+cr2ldQ0RfvmwfCVraIkKq7bwaVPj8FHdBDV
z7bRd9TePpArmL8mMNSNTB4Qu4MEbb1+geUWjveY9MFtYUFPmH9ni+tdkPepUW6Shr3JChzz48mg
R4ABOYtCEtV2Z0CN8bvwtMIByyIZVN8BXR4YGjzneWZK8So3v4r9EA3D4U/2cAkD7Hd2n2lRzBJQ
4fDcVGWidJEDZ5PzdZBJucmCGel+4NVN/F1w4W2KIbZuietKZM23FntJkdp5sOGfhzQi9KTNf2mE
aqNsPmAWoOObSIaFp5sLmWBl4gfO47AGwIuc6UlBTPCMuluj4WwCSspxiIrXyP+tBOZ/2uDkCNwd
VDAvFAA18IT8lILvJuBE/teeSuk6KSpQVPBKDiECn2oec5w+1hMEtDy8HNTQeOXGsEXRiUmsKGTG
MRs2XB4jExXsP23io0kDhaSSZgjJB2rLF1cgEsSWrOQn+LKojhlVQ3jtgQZyZwXOS9laRh2UtDqU
7u0UqVBYfPvvhyjdCnXghBFXn2MFseOdjquFQDofqQbNYsZ636dh5Vx1povX37pIUq4LYPNNClmx
ozGrQe9r4CZyG38M7qNTiNs6XusivCMd6FPzloJf4ATL+gyLNQUn5LsVc4ZzmfROlh/O6knBj8Ap
fO4HQO+9d7V4MUn3SaDSAFh5Fu041EJp6pr6aq7zKZ5uL6l8r1e8BZzTfQSK9WAund/eCgLcTe60
z5ZnhI70bzMRSSMcd6BHjhmC8Yotl/Ygjpuw7bnMf1kmeorVajg1aQLM5NYiBbDR2pfvwRNTL0cV
1hxg9hn/7be8UmdvWLdLrUze2Js6mAAjaVBozDnH7XW5F3/+9BLXCaq9bVGySHEXL1q2wYfgYPTb
C1RILpJUemYNVryoGndqbVo29PIRGz06kwwm7YSK0+2YjexZO8MULPNTRLI2bsd50VafHHVbIAlU
a6cA1RhyCg5a+TRgEqdwNZPRMAr/78cglBiFt8u89doaDMAAH1xzMyKSQKZpYQWmeNNPiUlarM0o
zK5HN0IKylW1VHqzJuvb3aDdZudw50EBkUNsyULr3nGhihDL+PCqzYFC07MFezU3IgmczlZS9m7V
XZ3ego6LD06SVBZf4mC/QnSs+FeaOoXEXYIgiLRngQNErkigsSOQAwwgKlKYNjaqjSu4OdNWuRZ+
FDyETtgL2ZhBEZGiJUt3FrBOPUOYqdOsJ/er4ZGjT4UwVDLeJR2P7uoaZ/NdgnN5ZF8NopworSK3
lHofseY2RdX8FT685AKeiwjymV1Ehdt6VPtjHjKHY9pSa/IBb0WVRePfszWr+UBxORoSNDoemhQW
toVqK3Mw3LRm6JrvvvE/DPwIJWvGZqnA/tRkYplDF1todtVLC8CNAF67ESqszMfMGarspuTLuNQI
p+ilOjqxpbIVJHMxln0FGCYqoxx0pPEyb6G+XqpZgbcbcQ7UKsrJtw0EkNT09x74mOCqmt9Z3dls
+BfbElq9jtRoSLhZjPkpw57TFeAMsDTczELrkk9kfy09+BMs9SE/f56Nowi3/5AYNG/DtBszWuXz
VZ7HdJmfUDwgbAHFrfU/P/NvOmra6vs08cYpLBgviBsEObIcrh7rxz3HxEBHvreiZ3HAKshd/6Ti
KWGESaFZC1gMoeWF81xphnVkQZJPlu2zl1Hbk3lmocWJYLNN2AxbL5yLCpcPGfYHmUg9SD/F8IVB
iXHxixcezQfzu/nkdIetcIJzh/7WOpIclmY4zCtdKvsd3SXXpJTAgNUAa4I9zLUGL7Kd+BT1mhT3
T1mhtrg0ZRkWsYrxhx8euu4yAx3A8vYrvAq+FgfiGPmAxu+ek4Bpkl4aqzUJG2HhwNXZ9piTa83p
a8/78Uwui6Fd/KTAVEEE+LIfN0P5FXsbYB9kqy/t9bcaAFEOqWUWe03m0zpq3HQfgFhrLlTCisMm
VIRkljp4KN1xgKjPfDaZ9ETCvZdWa++wfGA09pC5rBP/c0VWIgfhj32LuXEb6rtpOgiqVo6AzSx2
KKxl6qX23flmnKFWL8mD36ixaBJ2+BnRgY9pVSqaHTrRPANT6eiIvUYjmeYNPhABIhLZAYmoMKxv
1F0vmfskAiPsIkZqvrppC7xDDoz/LdatdOAvLPc0IzQevkHb4sIHaj4UzPEs7Qhi2tc066YTVl9G
s+LLhKD2k2pdARcI/dhRHlEaLVHwCGnYrRfVNNSQ95bKSmMY2b4dsmXc7OkR1mw7d4W3iK8jH85P
8wIjkJ/FEW5x5JoDfyHjZp54PQrcVt2CLTYcoCdOk90rjHlvvnjbiTS2v3rF5ZCMce+oZb6Vy+p4
Yq9W6M4fvMgiHGI4eHtIuLYWyOP+zh6iu0UMxhsnpn8WBClQQSA5XFBcLShJpWGut9ucCDgohc6n
sLRaKWQmY0ZYawbiHFCAla43bwcTviyVfMJtfA0XpQS3TG14mtgVpooo10adGXZtXaZz+8HYqjI5
vvyzA6A1qrlhq9t6ACkw2ohCmf8QeUKa3/gkK4ESBySiG+7b7dgYCfQ5XMzF+eTYGCR29JqodjWn
HCyHNjchoL+d/Eo54epO6vormndWVrwf3weBibCCVCHziz0upsEVxa0rdh0b5PtefCMRj67e77IT
NJXHaTuYusD4SdIg4kLGlk6G752KNnfKnAVyWFAd9aze/SBZvZW9/Umu2JE6c9M3vZC5c4BfOsto
lzRqNweqfAzm00Gz28hNVyXSFyQhxpJz/vn806Gqfpnpai4hOanZA6lXXRF41dU8/gsE8KFhWWjD
/Zjr6jmAL5dphZlXzkYzZoxL2Ll/I0OXrQLRJBJdKz8qt6xl8bLzmeWZuC2EjKhOuMH3BQcSdUq3
TaPcUf+FyovhwZQRFL6/Jn0+4OPv4kYUNkEzDKDiD4KdpQJbYNuwpXnEV2kW/4y/XfPWj6Go+KSi
QOd44s47DcL+Y0yc9S3AMPPzS6d6b2z6pBtaDZSHcStyYjTm000CD/oEcbeniAI4rAia+MwdWhLj
7ze+NTH6fsknfIsK4aFyls7FMtcZJyHSgsNjq2ML0j9eHrLNWQXjNiMfOGz0s4F+AFE+jgKNiRF8
DFAQX45c0TFKq3h0CQuKJu7SGNuX9jIhAtFy/cTNe8NuOoOYVi4B6fSaVvaLjuUXmBwOu9551223
GeUVdoviuj6M7HJ06ls8i2IYW4aN8XXvPzbvdOLUDmie2Cn8ea9nALYTmqsYVhjhm7+Ukg4f8VH9
7XrcVnDugV/lm2h9O7D/KlAlRrvGJHOSCT2isUkI2D6sZHHrNRD7GkwOC3XyiHlx4fviNLgC2Zgm
520ZRsSGwcHmUgv7y4Ynvs6vSJaQH5xP6hsukUKWW9NAfm+ubOVjaTV+zjzP6TT9GNHQT8hX+FTR
PvnZzuiGNjMSvnfC4OSGAMi2iqwem/Jhz16V3qSjBBSI6jGXnrwHGqxyJff6EevfMDucHBl88l9o
ia/p3o0fVZPwQCKGepLRt87VI63mWJVoN4o1kR0bXzGDFhRRYH8NqxvN8SmPM7bwHez4xggUOpJn
t0OzNAGU4V5h2HkaYoXcdp1zf6MNAQpqf/RshhhQbVneGeUUxRx8kwe281ircqZ/k/Qlxc6i8GNL
rZGjnkdNV4QvqKneAO03+2etsQmP8qJ3wVII9x+uCc+emO4r1XAo6IqJpxEDaZPhfkeuRy0/oPOb
Lt3ZOnG/kIgtlRqqDDQ722kYE058tRMm1qkV6y6nDp4yKGfT+hzMQvyGNr317pt2dnDBCv4fXjPM
vpIQpycuu/RRqdQd6YHJjPtd3bQPggyrPjhlLKHxfxeW5QbF/UcPnz0n47FlRTIPfOR7OYrvUugn
l0GUF+T0yYFRfQlMh6QV69eOixQzs9xHXuXu0jaGOvruYFswl+A9ImuzJi1D9P8Wo66IqMsxgRKO
iSq94cq5+QUnrhX5FonitfW9EsUAW1N1WfRGi3fxKvDwESpF1I1o/5Jiw3PksoDvGDIbmnUBoSdy
S+89GiWLuOhEKihGof7N9H29oMTBDx6l/rS35VGIzROoRbLp5BkTnvCrqoodEoPVm3n/hcd3kWrT
yiSxPG9E4RuzHQGQrPxv6/hyBAQprzrwB8v1l/fUd7KIZS+a6Ft692ecZW0R5Wtf+0UdNeH3VDf/
9XH1uTYOuq5fDQ6UI9dkQYlblBOCSrZm7oreu8yZew7fKo1jnKVPZAvUUWsK61T3qVACcv2riuyp
wi7KcGaUuypSRw9nkx9RcaT1TRZaXvML7nePb//gIJhOpybAcy96qujUpuAQox8inul0HlV6d1sM
Bch8lkPsACX/XMDzqd1ytiyFL/tlj10y8nEYJykcUgpos0InarfQmGNiQtgPgObawudc83PqSH9D
xMk0ZXo80tHIsBiXmmk+qFR/q8LJozshAmtPA9W8jaJoPuMGO20ia1UZf2B8YAyyi4D742hmVn+9
5444coMZZDnzoY3TIwv+gKNOyKi6ycVr9QwqQjsqcl3VSwqGkkCDWok/ICSarGhq74lWvQ+Gb7t8
y/LkANAJ+6Z7B6kp3eRHa8xcyMaVX3EGtnyvEFjiwJvwGQHbRHUcyJb47t44P/lIlvGdblV4Axd9
OlMaj9T2GLQg59Qnwgm15j+8ORF3rWBRNgacQXvFoycCqDVj6NhI45s69xLE1ngyR+DiqqmBQvwt
dYxeNq4NjREPYLtJYErVwF273XqiPninlDphKwTvFcEBOTd3BLlF3qM+/qTsbBWooEnpTFOZBpMK
fQoJp13gzOrbHAQ9G0PN3TYyYSQkXQ+i/CDx2TA9exmFX05JaW83e9oZ81NvZJJqA4GbTg3Lspbw
Ms11z+adjrwSzewOpFrI6doRmElHzU8rhTHOVG7+yMAZNCwxj/0U/GbYVTsjCHZcATMAhRtuBpXz
p/iUY1Gvz6ZSMn0+VJpfUnigjM+cy+vW3//AlUSexswtVfLKpVJP7dm8oDSBRj3/RBMv/UtVr9qh
4zwPwioc6eGIcpzxmPP1yzFmyrHv2uxSNiicgiWMyH7urY3X6HazfXHSZE45cTlcChFttiZfgAui
wZKf3IFEp3pIH218YdcHKYguIICOEEbEs1LHXFDSlMNMr43FH/TYIgc8Y8BCR4sgzbY/xR64Pz+d
98gSY97RQ+8gievF7ucGGzl6kbbhqnr0Aieu6qKdwcS4DKHe+ZfM4rUXfroCsNW/jSkCbH3IuAk8
2k6nLC9Wj5WOKtyYSNThwcD/s+e32j6GjkhhEYKJ/5qdZXcMk/zIGcsGQ3peSxeFNEXjzx3zl14B
Xf2J/Kt6OtQ4rM7QXgXMEzC8N6ccnu2HFp4bu27jGv+GlAsP1dKfPQsWP3ZGRX27HgJTwdfA+L0m
LgHfRmWBC2Yqr5txIBr+c9Us376pnCEPq4ZJO/cDMUcbZsDxk8Y5J/mbcM4ljdm0SaKcS4617U0/
YS5ibVT6tRT8UJiNtwSaKTTeiN4kx6UTQPdDPsVdnl5iEccWsZ1DQ/l8FhCOjulIvow1tJSZsgmf
MLITp/GXcueujrssaHvP2qD93j7lr8ZEZfn6iQekPJPNFYi1Or4OaKH1QgBoKyAlljwmF9qePdFl
v5WqKLtP9dbScDnkQHyTY27Z4Q8d1CFw28su+Fy4zXidqISGM59+bQy6zDDZ9bCD5Az5pdMC87MK
HUtfg8A4OJDMf13nixrnDm/GpVb1E6h9PgUMPlZKbwo2cgwkurn7Mpta5DQfSCATIze8I8NmikK4
ddDTb8T1Iuwoo15E4FoA362RafOL0jL15ldTjw1Gb4DtgHs0fazhOqEcXmSO8F27B+HZ1tPEGLCs
Srcuv9wlr+o4HX6QT+SRnSFLIBsuvf9Mf+cYRbS5VFaei6pdYzpkX8prg5XfwLwddJKvozzobpGI
SVwq/6xfpE+WnqTfY29b2b2R8zeJKSroQzChvThEDAOp+pb6Y3szY1q1UnPuMBzcWbRuOfE8/swv
fU1rEZv6Jm+aEbJ9TYT49eUziU7IByQ3J/Yl4rIVp7WS6/HgtXwS92Uim+MiRSPk5wzF2WOK7jMN
2mowEsv9/LWk4hYhnAZfXWajMb8kHlCSzGi1JqSCFviMFLwHRkZDkxu3zwpiHGiUdPEzO0QNlJBk
dy/6OiTxxvIExV/bnTx9wFlkVn34oI2KVcF7gVEkAknivwNNjw/O+MvTnxRdjJ8vL51dTsp4f5a4
Qla/R/H9RWBjpM8YesSRfwpjd7nGrMXVyYhQhD0lX273VwN2LSprgsVWpdCY3JMj3A0w6ieLgceP
wxEVjYrt15DcWLFE2eaxCH9qM7LZYUS5MqqE6+ggZB4A/90W/fwS0dRVqeTCEfSCVZpd6PChUxHw
LrB0w/SLM5k6h2Q536tYVSjAC82pq0SN0WAQscRzxXVcXF+Wbpm8TaJqHSJxPOoVjnGJbIwZRrMa
aPFSQ0v9SFP/UT897b9RKFsXJkCWxwDKoS1DyAfToOWttWr/STBXM7IYjy+T7h2eeQ7hNAEOJMFb
Sdymeu9RjHtvnIuYWBpYsSboZuwzUWYap9xRc0QPT6gsdWJmvGfQ+/ufePwCtJHka3ksY08szLDa
pIRFp1MoBn0uxsOAIBvZDoVYJwinEuSMyvq1O34zMijNdZfH9E+y/YWANJC/GFAVW7zZZBogzaHa
Bhxuh+/gqxNIO0G0wrcTxWTu6X11aXWzaLiR6AVCg286Z6T/SfMZ+rJ32k7uz5yxD/vIkzkUWLFK
MquUPE8PA+rfLh8/WymXabjYyiqes0eGU5/zzc5vjljWJEuUu46Irv7/BUpklXZi+TJZup8HVpiv
Qk7XjmcRYclldEMSimjvItt68qt+ho7CVcIosNaRI3V6YStxQpZZIlRqRJccSAAsqg6YewcG0FDK
vUeWdWUeJnFTb4h9Fx8QU2TWPP18G16TEjMp0qAkPIcpZR5ixbcMQmGtpJyd5OUmFW7NJuCfBy0R
R0/pkibGmWLQnZrhpTlaFcirA4vucJQzyBpynlUusMELcGtVMdXJRmhgy/mRfR8wY2YTyLRNE3De
xo0/xEugzvNgrbrk9Ml81Ciez7ty+0NW+lAcybaQgVRkoObZ3KdTc9LzHktIA9MgYOfHd1b7hAg5
T4UVoZF24DsD0LBbaf61M63J9lzgXT3lkJjP/XSX0D2kOXA2mDwRKEm++MuDGow6zZLw2MqUPXzt
piLHdBfg1fuVZcOh6hZZATn+vxUBnjnIzBp9LrlS+hRL5mLHcRl7JFgzgPFdnwB6jG+yKxV3OtJ5
jUkYw3b9kKm3HdL5O+lzfSW3MBDAytXZeSBXFG53svOzBvpL0X/jWmG5EO6ERfLn8q93K/zZIdJP
7smhDp0NeXL2bec74tASnECjeDHxD6ALeFicCv067lOulOtSnYu/5NNGrMR+/5hKP2dUmw3rXZv1
L0JjHRJOsFpDLitog/7LVD2wEtUhXtmUFOhdNsHfDU2dm2mFGFgCHzcFNhIWOvF/RKkV8PU4cfqd
cCCsab8C9LAjOYkSxus50GszRcfnxLGWRudxxRUVz7oTzmTxGrw/eKS5H4fh+rxVVsc6wPxi56nt
ZwaGsNNUS3ebxO3neB8YKwYA4j2SIMEzdIdQTbK4haxwa5xdjBFVlCD31awATW3EeN/m2J7WiVfu
9WfmijtlqmY0YowZulwU36HryXeWf7aEwVYRtE0XBU0iH9ZybYWtInuLI17CEDidJ/p+jZlggb1U
WA7IC/aanqld1jZkTbA8n+1ng8wcrpJqYu06yox3At1mz0/BVIYiy7hRCqg7gVW+5Romi0MjStvs
ovColyoh194XkGw0G19SImGLZyl1EXAxow7Nmat/J5OD/cjOgi5sT8u67bQeefqZVLydzuxYM+5v
JiRd0ui0GB0mQeQO2doM5Ysm6Ljgf+1DvAmGHSpHNe/QQmPyU+QlagzLJl6tJoqH86C0HqVIAs43
tBkn7eqpKrMzNzgaRx9A8w1a0QnKcD3huVGnVIekD7NXs+bSWYabcUpMnCcKgadKCw6yprUggQxJ
hylOMvoYZUZrIt68NOUaVqniSpeul9cQm0AB89lYWRAXdKVztkWpxq9VZF9/zJbTAFpJfF2Q0zD4
F+CSH3Nap51eQhKKTb0IK1B0u5pVAz2rc1dTcvxTAepB8M8xLMfqOVItLrIhE3uNjwywr6MuBXX7
k7tK2nfS7s5jUAIfniSUvnWT/DpUHI788Ua7lofgX4CnBN1UPC/sh/yQpP+/qbyDOrjawJHthxZZ
EZLCrqnoOkvtLGaMuOvqajHLgxuNc5xgv6jNS1SgCP5Fg9mjSH6LyPoUPCjB/y24MoK8uo57llFm
uJmM6ePaLrXlZiqSIUZXP0y2R12soEt2gTtHgufIEngaCY/R0RXUuqzlBqeed7zlmpOlCm9l/T1p
nn66wkYAabMWp01vnrk7l3qhMsRYq2MpY68VxJkJlclsKRmYBiN6aJvJrDukZNq7XZ0Ltornt12N
W9T1dnZL6U9wOoSqHY2KJTc1Lj26RaJLHbunB8hd4oQBKLLJ8xiAYufdqaXJcanUsARDpf0E2Q9k
b9Xa6Z3hUvWPE934CH/XsqCIvnfueNsowJvR8jxEGK2t7E893K/dQBSE4tJJVTaDrWn2c/q6s4el
31RRakQOGHimAA11+gGcQ41/jIlXTlB/EY127msNh7QhrmInreUBC3e/5SumJcl9w2BJJmn6xF+g
0/dOohdnBGgqY6pfnpUGoLOLPQaz1FWSmjfsYT4zH/bkZ/w2VXFix7Ccci9OVqM2l21DGDmJQlvm
8jTU2EyaNef7nOyy1Q8MIarI3HWETz2dJBaq9Ksz6AYmnFB8qIoGBdjWAfjqcEMkZQYKvF1XPl6Z
jBrf9gqJo4B0J3WKWzGqdJUDVVfxo6PWlmqX363kk9NXuVVvSG7qc+GtDm/cvNSdIkrOMLIWyZr2
sj5GVoAJV9cTihmPd1yLiV/zUL0RoT2w5bWNynqMfpVir6EfUdfY+ArXbxBn03FF5cIhK4M4+K7W
i2ugff21j8C7nj1Se2j+9MZ9y8+qUDGC0XXWqDFMw3z4xl+oTf9wizGvC/eVbh4V2MUOGjCLi3e/
FMeYBbkAvT/tq42IBktiiYEXbcTvL91cX+5Lzw6BtXoUKIwAGjzeyknTf1uO5oi2L/UomzF9cMYz
IZ3l3uqOQNWv6e4pKHjrxCCAz3erg7aDreMWdaZnJFjKNbnGnEyczO5qGsjVllz+0wcu2ZoetBJO
1lfa4RwOlaTZb60iyIENhZtXCKl9z/CCOI0t2pxQSeut4Vw+7308QUtJkIJfUAWAokctYeib5dvr
HkLmTdjrExqnYnPMI1grKTMVA92G4foK+HnbdJTUnwRgb+CziddyZ5PjUWwxcsYgUqtXcIAdreiU
pgddHc3PJFh//tdpVF2ZefsCtnfmJ2X/TKqFfAOXBBGmegPaXCm+wzVfHyIA/vvTsgAge834ExZQ
Kve7hNSKOHjqKKyjP0WDn5eSSdYcMNNV/4UcRDh20nVVNSEaWFQOt2akfU+/b4EzPmFEGH6gtr7H
xekgFF+K76KFOnJq4roOuG1oIS0Ysw8MX+7DnRguf0G0SEK4zKfqm4sGZOnyxwMoaeC9AttkWMdX
wuzHCxQfaQ04G/bsTdCr1xoIxWJdh9JuTewmuDG3/3oMTJEdcITAyqlSA0VbteonmWK88nZJciQw
e5b1B13nFDt9v0pgnqZAYknShVsqrxCmNUI9btK2O+Ih6oujt8xKO+la4QfrGOCb8v6x26tOZtsL
4bn+j6Gx5Ipeeb6Vp29nnvV1+wNDubETHwYsguDlVcMVgK/jLlo/2q0sggBi/Pd6OZ0gWuZBSQcc
ZgdB2UFmIB+iVC76g4eidoM1p/3YnTZbsAn6m+oAu24vlI6+whXJMhQ7RqjiZLJqqJlRhuKt+/tF
VNx72HW9Y4TyK//g2vn5YkXiQYoy63HFMYSB99IydGquB3KHO+T8r4hje1sGASgVTCLmkkN6SI0L
mVe9AvB6bUGaV3Gw7pmLh0S+rkvT1c+UvnwJsd1gwMKCV0mqT/aFnniBqwkwobF0w+6TbthnF1L3
54Jsz/IuLPSgEJpJp8e3gwd/LnxkL2+HxOSfJsX2PyMoLCbPxBk7i9XxaLMnofQaCLesHo+iMH5B
r+Kji2b9Y2PdxnzteYNIQW0d7kZ0sZ6GcZIOerilX85mnJ8UvkUD2Dfeq4eDMvnPsuvO4zSBMmWu
nGJ1ZQVgjEDWrjV9v/96Gln1jVvl5vHFOFgzQ30DYZ+RavUlYMuXsYbS4T0XNOD7nxY0QrGSsI3Q
5ScNxwK0d4eX+4A2GVfH45Qp9DoRpeqQLxU9MM1pWo9URcpO0uFOUXBKCGkc+xUeCQw+BItsJiqI
htlr/gT3Hvpi2IIf6XDFdr5BhWB6QDdNxjC/Qe/2Ebis9w3HpbD0+IeJ5+4KelluRWoy7sCifKFE
mIBnFHWqGPw5tJG7269HG3q94TPPjoohNJ6nsBobpFc1d6z5mfZ3kvvF/7vlovveWMNnX1vPStrJ
4v4pJZhgLoll10zxCYYhwLVhvnRfq2lolTxNSFhcrWJIGWQLq1U6nPNclFU3LaGsbbtIxshRv58c
C4jMKrbLDa/2M4ibY01p9O0iUf7IcnBoY9PRgTOEc8zFm2OEZgJV+Giz4LwrQTIPy3hH+pUjcwIq
/NOl5kXl8GV4S6UcOjpAsYkJerhhyu8WfNjbN0DsUcru1QSYawdx1PLlOGIyv0sbgJqrdlrJ3YJr
5tj372AsiET/0D7RwREXwV2GaQnY+v8EKQ2UcluWi+ltJWgVgzwenPxM2lg119DxfIMgM2QViZTl
M5HXWuVgYgNKQwZBUfy7gc9Au8Xt0Qd3THGzptdZI9A7RmRj1uR4FgcoR5ByrDcNGwHLu+olj/3l
g73q3YN5PSEnYuEdQjVBIBGqfqd6Oh3tQ6RHLm5j0GI5Ivska6NKWaa5SV4VDI14ztO+N/WeU7Ay
kSw3RH1sp+YgvGdbZ4uUlkTVjJdmvQweqmT75/k0W9UX5g+QOiVEfTXUVZLeYlpsqqdx8Stqdu7v
d+3Ui2MdFxxKfdTtM5vlsN9LTitGMviY5mvhMO9x9GJUZeEzGuT+WmXWw7cd34EVMvPYPKA2a8ka
J09YLGcycz2PsoY3nGwSkkn1Sm4T/uABbrtYi25PHcKJcdZR6TpYF3zFnSVGDH//g+O2v7kWqVdu
0s085AkELgO4kfZvdc0nnu5oz52MaysuKn6nVO9fIQP4tBIEgZekQqnh8nYFsSivCPTbsWc1FKiO
kzfzYMn3ZBcTE0W++wiYjvpsVJPwTcma2v5rskLJ1+2/GdqJdOv7MIB4i0ypcpiwhjsmwUNB2exs
xT5hzhKNASvjbhR0FX8tiwZ26f77JQnkJOo2TxPwwsVT8z6gscjI8E/L/G0FErkApnX+cULAvsEP
fz2vaUERxvU8bxBgUKsPdfWuC8WxJBknVue8xtbGzoycKW1sz0Wbm1qCcg3wmMNP8Yw6Q1OGYFcC
k/WQNSGOxnIdHaQSXaFJZXRJoSQKPBKj9OzHR/9UILtjoPsJ0xlecZsxARpFQQ9JdMGvjUB47tIA
PgX4oPb4gMt66FytRHxPcPJhEwsRTKDmHlZrc4VIAUxQ0ekgT7pd/2h2gxNLd07+MsyE7fmHMTZU
eJtddEfEAbicrhT1UARorI1ytrwxnV2NYV8OdS41eRlBDtvUapywRDRM3cDJZ4F/wx+rCZ5N/Lkk
xIlkb+NiHumAg65KPJzNAdImDoDGIIVaHA87yNYBOc0mgUwm8o1mXdfrMKOPV8iBihFjzkIZs9W9
xt5EfkfZLL9VazBO3nY/bp2vZOh0Zu0ENPB9CGvQLlW1NTUZR3LsGiK4EaekGiSZAtfr08nvyDge
FUAsCis1H698kyG7aglL3mtRF63ttI/qswFZvXdRbKawqizf5d+cGxEaRfGkXXQHLmCWdIBe/qts
Bz8fRM0fI89xfvpP0XbtwsItnJnfWfKm806ZsXy95TnwCj6TJs43aQ07nM7I1CrkBE8IdUM81w8c
XucN5zV7hOHHv597Ne7zOK7JiZKRRqvYlfec285FYWKO5+JJ660ArnBfm2qPXFLG9mXqMQIPtHJp
oD6j+xJSVgdaqMWalv+0qjFzi3HuWI1a5+qhPKRg8DmEqD5asPSFuMqa9Da/zSXIyVuocg5tddt/
Q6CTLBFtopqIhYAQpq5/j35/l3jEfsgoqL2O9W1R/RECZRDv+V90VVk2YDuUIsjjmP0SmFC23oGt
SfL4it/do9ZPy5KDEQO/JP0bYexu94MsQ6d9qqF6vNWfTuQaEjr7kGfukHW1lpSTrRFYg7G+rJJD
chjWwwuIUxGwSVJDLZhYgwcmpOTL7qmAKfIxxCyFHYAD1N1qGPpdM6CvkxIb/WGGYwtCgsl60n37
Tq6OuTBly+IZFQFnmBQj0unf5hjJ8b7SIAOpz6Zp3pImOOK+UG09bnF2sWo7CW4hGntf2yJlmUv6
V8qbYngrjNdaCCmzbuEO0nGcvxZYoDNgJam8a02cqWQ+/bj4B4AkDMgLFMIVJZ5brryJDLHcQt72
NCBKV3j6IFSNqtogcAsHq06smi3+TZiVhCmxeHutq02s1toCC4IT/l7qovZpmy4oD2Z0VffRc4y4
q8sVMX5OJVyEaY+l9rb19HnVkuiKSRQMRbhHsyvIxo34xqDk9/LzYqxeiReniAHEKrO8Srvh0CgK
+xtJ0ypme6FwfX28miSeF/6jw1psJPJ4AcquAbA3bV4weXflZj6yNKrlVRz26uc0fdmo0qHINnYz
men8NGTl7Wmc0BYLcvJW+GEQpQGGJCV9MJU9+ctnZgH0ZBHmn7ZjKRzHRx0E54dyYfxGAsfD7bHH
E93uTyk88LeNy91XH4DO5yYGI+g76spDWlniZjoIgyJ/M6GqJyNil7mlxuXhyPv2MuCWLv/3DaE2
e/VQGm1w1tCSjorEA4AFZFGyQ5/uJqB5WHDMIPnMHLw/tVsBJZ8JJuDjv6lckHqAkixe+z7llMJF
79op8QAtLo5PfM4b340UVijY0rTAhpN29NnWuBIZHigzF0M/j+a33fjsNClse/YH2oWO4C6tz8P1
KY/R76vNTdJdhc07SyxTopvOqb2bbbhUAPNTmYWPsr6zHA6jFS46O7qco8LKaDIl2FJWVGsw4Elo
ETYUrfUKYjx1PNfn8oHZAD7XLeRmHu+ksTuoB3Q0jGdz4tgdumYPh8YiILLZJuB913TB5qQ3h9wp
v6vUjlXll6HA1RZQ7oxCSN8f/AcN412FacHYOW6BmWW7q2mygK5iRc6Uxp6lHyHXGoorSWvVcXqq
E+ggIgfmgBAdT0GQ9ccxi972jc3jMEMvkIDS/N5csvwcOYAo8WoO63SSau6QHyxwrQmd2Q5WH78t
o6VmMMzCkXQRjhtpHSu1jilDIQKt1KAkQ2EPAOk7QC1s8rUCxuoMYn+OJ851Noi59BTaRP0WWT4w
eFKikeyfBsK+14XL6UukJQZLvjIK/C23CGUQayDgvbltOkPjwnNy93pAXXv1GJ3tpKEg6WQZdhb/
Nh2p79bUCx4e93fksMXHUGcr91FdmLzVQqJo6gRlHUnZqnEFO7Ry1Ao8VfDTblaFGbuHEBh7t/nT
srd183G6Sfmx8aZvk4+veaS8Zgp4GRt4SgfbfZwq/cU1f9AF7SRQ2JTBvQVFg1KozOMY4/rmjmoX
/S+pBK8V7KKy2ts+ArsNYpMPJy9pxBJPJvHtSPP15cnlaFjDi+MCnaRs6IUFL3ePAEtiN84LZm9f
FMaYH8YjzBYe2PdfTkA8hSmUV1NbkLEKZnG1f9UVBVJjL/gSU+BjteDwlM75MQ9Z/o0klXmHxoM2
az+n7u133QKwp+ulWTUF+Zpgqt3Griv6ClDLpHXzmzn96ukpwkzTGruHVwOyUzcRaLw/f2ZoQt6y
Y5mB+5FvPMI0frJ4ni1sA1aRem87kMy8AKFRop2rr1KqCLJrrvII6h96zh62C2nsv3XT3XCZ3n3n
lIMrpxNXc6RVmeFigPIQZjexCSYUQYkguPA/E8vvj1unJYvNUJW5ANbDYWIKADEHDS4VsImMtejL
SV92WCDJozXfSBfs8rtWmXRlfqXCl4r2NV4JmqjUaUf1MjFyGhXOqS168AkfgCLJsflbKpLVzmG9
uV61J1Rqf8AYm2OWujoilk+yvklt59735yPvDP8jj3Sa1x8i4OPRW8HxBfMcpCZs6UPbNvrw/PdE
TGpvlIzFE/dZL8C6+n/ULfma6MmChgpQaHLEUaAmq9mCAmWOVTw79yfroMA/+2RoXNYoG7FdL/Qp
cMdCSyU+IATGvq8LOihGughfmYp/YN+oKI7KUI0cJWRTeTx84FhXoUPDFYX+/Q3i4kYTWx8=
`protect end_protected
