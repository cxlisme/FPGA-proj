`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mPx7gcQWvUiXAIlptcS0ga/HwxoglSwZPSAvh1Lja87QFX6EO1tvAtW3BEg2Vp3HivYkp2SQvnX/
wf5IwSVugg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
u4kYBbKWjVmoqUxGQIVLXWFveYVGjS8KXANLcMWW+aY7ihS2tZxXnk3ijjHseANEw/GD5bURIhkJ
wHNHgMafDMxk4PoyqdLtqxy3iP9j1MeEpH9OoyR56v6qcdr3P1DRazxtJ2ZaXaFvkJSsMWBDAVQb
EAvsPUwG/uWyf8K9wIc=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rcZYcqDcW2nDRCEfMQVN/Fk1OfFW875uC6ei3MlaCqhRnkhzT3xNk2eZbf+e+AP9hFcz4gOesi0n
ZoKrSwPNM4QWWQUwJVjaO8mmjT0knl5bHqmrP5PtUa8Ymb8JvpM2TW4eZK2Uprb6QEt4vqyh7TOP
vhbgM0gvOVsfurZr85pM+sdQTj4K2NKqCt95to1VCJH/hGDMuK47cP1uzcMQplSPzUkPukYqc5u1
65JQDYRjOTqX4AbM+yyfDWw+pb5SzcyHehsXCJH0dv97fYVSVVRFHixh5JYVGcKStfxKGzXXKQhy
T709LnMhsbkT9A3rMvt5la92JFzNANaCQ4q3CQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g2wR7vfvAF0uDhoyjP4PFNh7OLccqK1GsJSoBjOisux//jU2ZxVmLxA1YJAl8lw4jONkagbbp+bD
DeKzRS2ZhyX8p2HqWKvZmJlJpU91NNfgEUeagxdfB5g/ozhVOyy8QGxIiIMb6WrYXhYmtrxZNloB
n9TcaPYLMM7L3bin109TK04mlunQYKeEo5HzUOQf5KJ/sqzhE+gaF5v9vGZc+iE5PyzEZmTRiFkB
DIKvHD3bWL6nrSBv4kJGEMbH66PqN/cEKc8g6Vp6Q1KwRoVPABYLyvfgScY5ycPGYtzU/pyN140X
1iUlGE8ESrGXM/xbywed16jF2DlyQ3LUN34B7Q==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QhX3pm1tgaFGdr2rg1UW3M/brT66TBguCgts2VP6sg+tkLIps/ZujQpBhLiiUBuZpY7LYUF6Ttcq
FSLxzJjaRAKHhwz8QfNP1LvV8beGlrmElSBg4WQ1vh7an1NBCIV9vJQ12Jb8lKj8kV4h1jtFHmSH
K9jxpumxvGxg8OkyiZFRMV7wxy5Vgb+iLbXznLPN1sO5bxy9oPYkEE6q3W2XOv/+6RQT7jrgsgij
Ryn6WmRS1JEb//SBh2n6mIErQ3VXcu4P5ctFXtDE8hGFBRyM1uhm92HrFtwOxkQS4cyQYHYO9iFQ
G1fTJnB7JigyDvGKfvwHOOMtLjFExIGVquRFGA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qAV9ax+P5GkwGl6RgX4q3QljQNwnp3qvuISp2RvaZBQjaPrHqbafHxa35DhyBrgca2jSUOtBUvJv
KqsgFgfZn9V1QbQ0RhuZfQ0A9iTYX/dan3GdDTQqO9dUx+ctLSRf+zGO6pzzUXyKS+BdkWX0VK7T
nlxUO8Eglcs41Aow9Bc=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ersNAxW2yyOqkd9D0cu/x1eK3Xnna2vZ+/lR7+n72DdUl9LOW14owvbVJOgkJzjQh9R7373dUheU
TJqG2Bj8ZCYCqOfOaa5QxsPGyvnovZkK5DNfXSZyOo52a3W+1/UREYKNJQXMoI7o0buPSR9vjzfT
VP6gcUF2vI61llqn4hGlzHjw/Hxc7DZ2qNeQE9EkKFRPZZAg3UFlr5FCYYM50n1xKXOPz1GiYZ1m
fQ6rbSyWQGBnCD37asaeCyMWyupLe9e2+ig34/lXawgR9PYogJ8Af3Xu1/jMBPPEu+9fRFMGdl/y
WGXnDPxDcFs1W3SQMXNmK4XHz49a94IR6/sTyg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 133280)
`protect data_block
maYCr+DoYRR9+e01DfbGe7eb9mpZk0inuCuHyigTo/r/m7zGJNWibckAOyig34fejLd5Ur+e5nuA
Pe5FaKE83SiBWlNig7YCchLQTn4w0MBYceCg89pRMV3Kzw46EpyblwAj0QVfwKbBJ+fFCZ6wm2hO
I8x+0dCk4gQWPuY2vEoLEXSbjHo3zSXNcWnClY7h518zzuxU4DKTfC2lDFNwHNyh1ADnaR/u6vLZ
6GxoX4oJWNi4juE2WgZjcgHiWkuk2V5lJGiZMpouubcE4e4tPwXSSEA9INzNLprTqTH9X2aJ9Z6N
Id5J8iZAarToxESrJBhSdw83q10gFPcdEXjyfKoGEpLfyxVxBC9Gn99j52Str4gT7EPNP7y07pzf
WBFwqAvZ6iOOMPIenBEHfnlm5pRZkPr+Nrv3ns46RdI2L7OB4OnZpSJolGNSncwrrwr8s3r3qbcD
BBSFEFqQgMZOD4OnHsJB+l/2Pp3RIWmImWA4gsHqGDrBxvlomWlBt0m2o2P16iSqTE6b64qC2ksf
cwSvz6/+vlYi9uZvZKfoSJuieesxkebRr5vK1ka5BeIfgRJQSsV3GT7ixyzgPruv8YlDbD+WwER+
3DQ4m9uuk7lh2tZdSQU7EdyAwDigInQdvRIBi5L0jSSvqWLb9Ic0ilq7xocoOKRsMxOcskKEB/NW
cei+1LQT2DrPqhESBtge8xWjl6c7Op+evvK7LNrhqFdLWwWl5Enyt6a7MBD2DG7hkCxTpPIBKMIK
VHSRkj3ERsrQoPZXWWeylh+Hp6C80WLPIyrWdmyb8XQszq/V6i2o6LrHJdyjQaprxIA7OonyyRlV
Jh37TK9b2Rl2eepC9C4/pMJdyJ79lOBTm8NlJZ6eSx7+HIYZiKcn3cjF08/Qyid8P6YzmuXRe7wX
1IL8UEnQGuNLnBx3A5rr3XUuemJZo61714goeImDyBoXRKuBw7veJisuFMyS4yW5nsbeno6YBf6w
+QwSwkTEpb9POCvzufzuvw4Y3QimrKiN06zHpJLXB8ooEVIb2q0Wj60qW/Qx66VfkjIjQXbjccqi
lPXj8aT5FjjV4Y+5ZMoRnspbCAc5R/XI3BFlBUkec6aZXepv8LGJQPOt1tTb7Ijv1GwqlBf9Imk9
4aKegwszAHesDGnFon3XkTp6W6BSe5DpICT0+UumXqWxG5UEyl667AmLZzK26ETrYjEHJ0GMT+kf
1yW1MUZOi/VQoAdQHh45QEvBQLD5RwLw09G4Oqf/9e7bCtooJakf4V0W/tWEZbmxVq1psW2SIH9M
xBxe8YV1fq22OEqRHiWmLbhhFL1VEp19sIa2sTpv/WAdPtrwTDymk8sP46DLoN9L5gNdlEG8/gHL
nzzQ9oTiV9kOiHd1hMWaYO4qSLuNUNHuOcpyUztq2bQuZcvzJWcHDjAmxZLZxgYvM4+KaaD7jlhK
Fyya/CFYot3sj6Geue9m4fFYZENtEgpMZU2XrVoef7Uo359J7WfuWP3acypo7KPJREGjVknirFgr
IYmSVrOsSf/lgrE8nX1c8Yq3yBv61Y94lcw92lF8KwOAJskqcqjGxCwRKKzh6i9cvRLEALb5fJyh
G+2C+akhYaV8vy92E8ADDsgH+/svwbwFvOOPSV8Mta9iO6kSIEyTNhGGekks6N4kAUq007v3Vl2J
NmcXc9Z5RxQvdWrDSJYwdtlzZfYQTMg5rQKK0jaOvIr5Rj7+0dcZ4L4t9KNPvsdZpMskxabDnlpO
m7+ZQFpk7nwQOJau4CtD9WxEq76IWMeo1UJxhYdAOU/5ADdBMgS6YxGR3Ticr7jCoyyUFCaYYrzA
qav2XGq7WRaJoFERLdZaTXzmBuGa1uVF11PJx+0B7HNJ0EFeiIyocEgeEgJNjcY3c+Yk2SgMyygL
4odxooE5f0UgkdOdTea7jxQiMGBv23dnb1yHiqViPGLFzo5oJCjqoEsBB2DsLbmBweUYQPyVc0WI
hJvUnZcnsU2fwfSulVgudasCJqzQzcU7P27vWZ0ynoxNDuo2JXi6gvwQS5AN+XpmVwzyo6/p7OwJ
yjpUThIgiLQ0oPWOhD+liHGHBR/RIlMZKpI7ORTYq4dOQ3QMxAcqKm+JCcN/QWIXk6UFjiLnbTn8
Px7kElval3GZn0EeaiwV7PjFC6MBkP0pi6j5OdR9HRNPTzWseaatwBPurKDWvK6nUsJ6M0MRHwqx
3zpIq+D3bpgITFs0+d4RAJjJG6wbpN6loRlPign3x8eFMBKfIAXUPYy+vxuyeem/7i7MFy4/0CFK
U93kl6ym9UJ7f7J0+AtQwWnH3Rz2g+aVpqo01dJLsXy7HhQywzOx4RzIeLEg5nCeT6rvfNZViuYl
LK+8skk405miUonw7UGCKmbJAiTdVECxK5eRHvskRalqOzA+XsFyr+qa2h70QPhJG5jqHRNbPqgB
w+pQunx2F/O3TShdABgLAfDxApZAlAFk7HdPQc6NyAxhlaPl0dToPtqLuqXi2qh4d/6JrVOHciqF
8E+1vp5FlFtPCF5Qmx2Bdbybqjxe1y9614SayuMBzuj/Hgo3AEr0aSFGPvzxJUj1tIeIQchYhd0z
j5L2CtoyDZhUWU/0h6OaRY+tgSwof8BgpakS7mbP/kiO/3Qn16O4t/oB2fcFvJ2pyg9YBmx4cVFV
p/u2SDq2+p0kndM8srToeouVU1CQ/DhuCdi2iUnRcNniLLBim+UcChp4yVNe5rqOutdP+ff2r8Q1
TFxqgaADWEKrnkwd40oNhDTMXp2vxUzU/sdqYEpwk3bhfGcljCV0YvV5C32GA8ECuhy1o5OoKEXD
G+7qLuP7V216xqAzkPtuwGEhJm5cV+2FFizfL7GX7aowCLUqHkkPBCTFHOe9vcMCGHBItNeUKiEa
HMsYSyEyY73xdK2VYCq4RgvGUHvr8d08gUWZeS4iYQH/mUMuj6qYT8Og90Wd/KUdHpxRqnJE8/jV
duk/wVJ6xzYoSzN8zenc6lxwHGxrnMVr4c85aaP2HXvn7LiK1F7U1sZ9p50vtGPPVGe+l+r7d7Ht
+SevK7/ePUpVM5T5y9FV4H7vcoUhLIXeB44QQgXoNsflUdOrQftdVdpEFgtYgbwDI0h8iL3VeomG
P3siNzcoh9fiY9E5hOEHBiwJJImPilmASAIFozfuM6M7nK19epPj0JYQUIlq5uIZv3hYlQuIV8Uv
DgjjVhMil/OaLYplODerG09gHvDaj+tJMzBTOAM/zPzLk5y2DoE2m/ii6qqy3XpjHNpJnre9fEKR
W9pg1q6cJg5lpdMDp/Po2RDPrkBudbk0c+yzLlt9UiiLAI4WSqP09NNdv+GUUWsIwoqoUaXS8wfD
39QebiCCJVkeyb71vfYoFNGYNlqOTc9jYcoVZ4uKjU+lUNsQT4+46zdyFwMJoz0gIaUkzvmpsRjn
xtJdiFoe++Js3ylHivAV25ZmHLGhlEps93gOqHxYmP7SDo4KsrotPkJ6p2cJ6Sc6J6SMQBrHTKYs
JBupdHLTnjU/K3+azTTNDdwIs0XF4heomIgnQvI4KPtjs3dfWvWvJkq55LQLbFCW8ezcUbCG+kGK
Gya3LyHVhD7hlVPPZ80svIiyZPXiJE2w/MQq2aDpkzZoxwaH6i4qFxgkX/cZbP8wroWShdKI1+AS
edEolCJqcY8BGGnApKTXuMoeMEJCUMSI255fgFiXn/goXR+1LY/wpjzv0Y43FsaluWzxa+Xjj6qK
udaUzEaf3FywcW/wY2NOw8L4pq72eoF25HU9nBHyW+0/OJzqu3q7VdtVca9RRAqvF4RxY+JMgFOz
9FB275tgd6sLGYumSyzi39lvGgB1vaK/iCoXZru6XjacUc+KfLu2lZ9H+/hD/lpKYcUBYkQy/IMb
7xSd+xRNsl5a+RePMjHITkQN1ZiPQnyCosyO4kj2zy4jl64l/BIxhD3mjQYgiPbs4km2QRetZ3Vl
eLjd6RV7NtZ2Oh9DG4tMRNP0h5b/rdqQ7oUIPEIIoXRjR5xtkxg65Cnp41AVsc3yvp5gTU/VsAeg
kPhpt55sNBXgj4VZcj+XyecbFNMTZg6sLPZZbrNw0AvvOBfwsMwVCpyN9RS/eqKVq8q9hiB1q6ON
VZFe+UxQGQjroKzcmUFcCNDP7kMeWHKkOyz3HNqlJbHr12BM8aVGvNlHrb5VW3LRout9u8vPttb5
6TwO5ajIDKurzi8g+8nFS+v24lbRZ7GOVlObcl0g/8q+ZEHMamWdcIw9dW9sKc9il1EMfj8gh7Gf
keZ36ZJJlZz4z0WOQ8bsI/WHIG1RBf1jVkiQBAF8vSddYD7AN33Eols5eWbkAWFIEk6KuY4Ps4eF
7i96NJGGoVXQvK2fpiAcgaqCdPPuUDTw44ea861aJYlxGg0w4LFKerZfiR+gz1dz7Y0ak9n0tqTL
ExLNr/vWtnJ9uohrr5ulrTRJDNuTGwTGhauDGesmerw6l7C968t7NaeC/JbiPRjSunkyaMtMC0nu
mAco6e+saQlvqvIy60Sw3mU1ik6n9n3WQuJVX1pYwALAthGgBCjA6G5/vFFOuHrgPXv++aYXx/aP
c9lmkAzs5kfp2uI/+T8nIFFSkRrhCOLHjW3zg9muz3pvgf620EkrQFGjLoLMvG29Pez+LOjef3EO
WK/W7fF1PIa+QqiA9eZqs3I6OZwhewUiGjFgPMsqPqMmyK4Jhe0r7cgIojMG5WwD/95sQAL6vpU3
aMJsxnZLhb4k66Y6Ws9fwGGwcB2lBO1QJ56JzJmjzF1o2lvE6V9tNWEEP1TAamISmjkFEEixlhV/
+LdWyL3BR4fGtI3rX9Ix23oWvNOjyiUfd43jwbJKUngFmOtzvy1mvm5lu3Zlj6IFbDQihnM1GR9g
B6jRIWeHTYg9fF2yBkL/02idjssfplI8T0FEmi3lsnEIxTi6UM4c6qW0vEHuWYqRjS8IhX+ITHUG
rNPVIOSQD8ruUzCmGEN4/o8cXpsf/WUmHII4h3cIh0EXq86WrUpVcW26kX08BvYKWGDe4ft9v6P/
fpO8TADG9Le4Nuu/Nm+EhDhvbCyiHOaY3ePwkWL29N1Xhlpq1V+IUfqdQQcb8bylAqVOYFGrw4Ql
hui/tLE7xpkSJgBDnwV1kheKjaa8HFyWqryx3evPt6+i2j04OAZ280ivdw46OhNytfJ4oqtKk65d
OtEYSgWf5KTC8ZjNGg8yVtyeAK4aNA/2U3z+MnoF6fuG51+e1lAIyx7s1eM87aThJyn8AN2+nTx0
YUyGbh4OkBBhr4IkDxlo/wuqG/YvNLJYaGnJ/lUa4wS6ComA3++v4AfaGtQn/GegyxY79IPUmANZ
ZfXy4drJ8e5ZCho8L2DxwfBqvzPXXzx+2Sk9HX5cETzd/XGSjtkd0DCsfdJMasWLNItECZ2rn0In
tMp1HmnSNEcRFozr1kSOXPkVnVtMwXWReCP4CKyvEq2kqj1W9EAXAL0MzbnoQH9nBtCuWhi/ofEA
B/CCrqSQYCQWUXvSDX/YqpqLlXFWnF+6KK9FoX4OYEioNWrhJi1XAkBuv5jJZNpNgmX5MbbO2PAO
mcr+4uJRjpy2JEA4GpsaD3h9sYrpkmKeWSu4e6yNjiY766TCuYH4loUbUorKn9cKSqVhdgmftVI5
Vc8X3ErOLtEmbxN7+TUi7Eth6P7fX5rnEfx/AwArmmVs7tc+PrGrEqfX1jWJANsPGB2NPAm5bOdl
9zl0B14uTMAS6N9uY+k/D3+2FVvCkfupTrsIVPjB4yKdZ6vxocThFZNEss19uzyphT9LP5Wp0XMA
EgenpLm4NHNf2S6fbljyJo3vr2Cpd4kFGwyjH/hIex8eW5kdKNkQWU8o8IQtiFrJ4nla6uOcOy1G
WM2do94vUwuZf0Sc0rT3nPMz/kb6F5gfhtncCPzOxg2UhEIH1KVX7ln2ROBrEssqUOiJuhN5oJN2
Ig3AB0XhuLbug2kPwxqapagC2eSb7SKvlyusI0fRXBezvlXqC0xKfeup6jnL61G/adIOnTITWjTI
Regdj3Jo057sJ6eEEPIjN05xnLZyC59vK3rtJSgkoZQK8srps4k8AIhPRtSMuRDjHZqnnxh7VEZq
1C4abqgW9rfHsipU6lEk4nZ4xqX4EuZccmGNyp1j/hb7C/y/6u7dG+ImiteYySRbsR43bVoAVZw+
s2id8C5nY2TujpNDSm9oraWZarNTky+lY3SJ+6icG4I0t977Jg/S0uUE1egM1qD0UPQO5SQSt4Us
gHuI5NvJSnI+k8zvPUA8Dus56rgmEAsvyccQDlMv6wv1b1vscQSCPBV1pGevQjIzuMwpYOktQUqo
+6FgANbdCnJ+zDRE0AVb4XfWPMwTcD7GLn0TbKozqQ3/Bxwi6Q4Co8Im3NXdiBHG5JYCZ4SzJ+YE
vrKG9AwDUHBZ7j5XqSHYnuFcku5GkIUSbM+2OB8FmFpZ7WjAS9M5QjWo+f5PRuuHUfoXxLChj/9v
8wga5QJ/DidVNhD8Vxg7EXvQrFH4FkTSWDivV8n3PoeNdIp/8g81ZDUEV8KDvbgzxVdbVJf4KqNd
aObXKLXgexud1OQ/3n7IukVoqa+mhYah+yAl8LT4jyCDno6iabn2YHdYnSB4piVfCg0n8jVVwtX8
dl9udDz+wlVitUlE320TWDVRNJfnjHpNUAeFaCaVsDH6HMJFI3ucV1YEmhbSK4aQk481zj8WN9dy
HsedMUfhgyO1+1LoJlGofWRIzHJ/joexJjNY+ElpC0rlCd1k9wC5k+Qzat5rt1JBU2izh4u5z9bS
WM1L59WKzMy1Vr4M4iTFEBkcPMcQduljf6cOQV5IykilEzDqdpy26M1JJUDQ9+q67dPmzABnDuI+
13KnUr3pxiGIHbUh+u/lJYmxYQ9wfdiydjnOq8uobkmQHFaH/HoBYMzaP474OhcEcd7fL5yA3/wh
pl3Y6CiIB3/jeYnzUsywnWL2C7R/oxo+n+c9GvOMKrwU51jsoI7bK49zRFB3S1abpIEYP97vqFrw
qcHhgOvTwqEbhnn+ohVBl29+kk9ikSRRSYuySo3FIguqlrGTn160JxIOv5sUz+kkNLhKzCyGzCLh
fdFRNpvIxDY5YyqpKNtam5KkA1jhmQ+PuMIwVTvQXjudW3jCa/DCwsk+Q+cSu4kQR1zqw3g6RlBv
3Y6dKrVo6dLxM3QiiC4rM02L0diEP2KB/HbPypUR8n4Okxl9hMsTS3ywucHb7fdtjK6w3k33tvRv
BjtyXI81W/FIwnZDjLkmmxvkImrtKfDEMXbcuuHqN/lgEZPE+URwQwZijKrEw4VPxjQpYZDcmWuO
cpnTpwL59hlPL91g1TsAsiNWqvy3DWfemdI0mda51Dr967uJ3UmuSP1DM1JMqbPBc0i93r1dIKZb
vcR0r/FnGG5tKjiqIHTiPGQfLPYPIdiqCoaDB/vVPwGS2Ox2PSJc7vARsHwxNBzrrl/gsXPt+tuT
gV8LBqjJMSA/9mXkO+/iEvf/ip2hO88AtAHDIwDBvjdTc036Qlx6+9d0+NVQXOp1SDhT1HbxvmMQ
Nc4hIoEo58cIGXCcasbxuAoeS1hXQ+KNIQ/wMZwJKvySJzfPVGgtEX+HarWaI/tgoNf/qqri2Kgi
8Gioej2EtIxeermB/GvbAfqBy1LSObUg1Tm7gi7EQxNWqNAqQ7UgQ7PUVpOH6hh4apDjqoFZ9ocF
9y97AfnDYU3OBPHQAINxfQf976lBDK/v/GSOS1lfkNdLedWDMiNthtP/O3jcJREfYgPEydOF1+Hf
+UB5tRW9SIWK07ycz0vnBoRNzik8eUJBf6X5kdeFnvXsisGolz7ursaZD2/tSOxRiStcic/q3yOy
tw+AVhcPGYK4gm0SA6JOzj0PcuK4hUvsiAG9/05PSGD663evkgMl/iE8+VVVPTgwL6umAiaMuEB8
v/ZG6Kgxj6o1aiLnhiupUZkwPC1AbQY0Nq4oQ6Mv9B31FwdyFELNnK8KPctYO0djZMncltyApbuJ
UJHpEBAZBrR4cfqhpxjmS2NsQQrLwFnRzXgxwOT3tZPTQ1Iv5aoV8xjScayCUg94le84D0xz8iKb
VFrnHLo/YI647C7NRJzMoMcPFLrXZccforSQg2r4DBgU7sJMTMVeiki74K72H9uTLVqZfVDuSuQ8
ZC32UIf3A829MzhIPdf/l9zBksIn69HxT0sxDP3GRybu6zGRK3Ip17gzU19E4Q3gWNALoik8N4XM
Gtfv5WthBA/NUc12yjYPtQs+YsFtuRsRAYgYCSVNEab0zGgGBMcvX/3o4pK21WY3+i4974FwDwJC
MYiI3ycwOxnw9rMBcjhkmx74nh4W8OR6zoVQLxgLgKlRv+UH6M+uc4sc897kHcPBgMvlCPLphyRj
IqbPEPJ0y8HYsCe38/gq4y8txqaq88i+N/A17tEX0TvTTwBnVUbIUitgIMfaDtc+h8yJ9J4KuN3g
zXGl7g7XN9tAt+d3BC28vfQv5b6VdOmsa5vH1XCMitubKvqmu7RAO4GkkQhzKhr/S+REzhvi5CoF
3xX6ORn5UQEp6D7Q+v09ZQyeBmDNK6I8H/29I0Etpuj7RAUvJFL0gBBrXj1jkoP1wm1OYRkFx3vg
P0pN57Vmt0EsG44Za9MJtOiqlH/qAj7lCH5h+zijQNjdOU1ZxAI+y0n3w5+XNz0ALqTXmWi61IkH
v7ZWkfDwBKuv4mVC6ypjkVD7FEMKizoZvZT190frQbMyRZL799QqRbMFCdEkfuO+WRFNAc+BMwSQ
UnTj6Ie3Cn/nQ/eZxzvNWoauJ2GEbG6mzwKXTovnvalk+0mwivGCZW9mG4b5ewvguZK+teE+9EMI
+BCRfDA1roPiMwW+LRgwmeCfjTFhKZDrT3yuskLvDAkdgTVRCdmPYJph38qMNigVxteLePOeJNcC
HKzAbEgjUpzsFwHa7aQXd0RBOTdPuFSOI4ixcR/k4xv2hfwhT6SVcx5xjXej+otnFc4yjA+72uJp
qSOB73A3sqsOMZTl8FVVD8F2a4n+m+jKw74ognrkx79I/1IO5scD+qS1tu7RqkLmFvuA2oH0QzTU
Cs3yRLlAYmAf1P+qDT4oAM97WjQCa6amxiIUD0SHDJyMNZa9+96dNGENDQuE0jGKbXYjLDpIT2+z
UUbLYvkIivatExLgM55Zawv4VRzToZFFh3F01om10iTvBCqTh45hfExkLweoig55soQ/0GoWfvhN
novjQa64863QW0S6FhBdcu2dUKshrCW9GDo2/yJ7gz0gJrfTiF3yrO2oE5rnI08maLHTMIUeExff
hmqbsCaI+7WDc6pnZS0fb8+1o4EIz7yDrkxDkyUTI2sIpmGHZ88/WNNGW26WsHZ4Cu2q8le1UpA8
4QEtyjDppL1m/iw7hkyeQWKlblu/sJkk6+iSeFmDE3tig9A61TgQvrs6/jmUiC63Ue8V/x+kCLhr
BAJoWp1vrZkIlvkdd/UnoybEEQ1yKsBjKaZEvV5kcFuzXWL5z3UU+9/2yBKF68gqXw+zzNHaBuZn
WNkCkvcRbHHTZTPF+yUwj70noMtkQa+Ysj+AkWvDuCywuJjccnAjeGXpth6pZ8naVoe3o1A+fxqr
TAfiRITjeL/uulhBPagQSEkRH1GvHANVovIup55JGTVXOQDhu2K6GXl4aeK7n8w4NLbS3FGgwvg8
rz1mEGdvyfVsJLo/f7VZfckPJx+46pu20bpFNWRGjee17XURqcaJ0qJgVhWjg6awsy14uusnfIXZ
tmAPuQNpSeVhRrCLeDKx++DFL7ixNtb805P6Do6nK2YhTJj/QhrhiIrzA5JfXYM9HSs7MB6975xR
LDL5+QU3S7EhFdPBLgMQwLBbu2HQFj5U5EBbtRWb0k23wH7JXVtWu4Dl4Hx+4BLuuSObgeJY7vWZ
U+wF9ROWZEwyd0HIXND26IbBmYhCvCZnIh0/JiDwA6m68yHzpShgS8BzE3QBt0fk++flmm4qxPn/
t4usnFEr+d1wq8J5O/OPs9/XIysHIRfzlF/C00WEayU+qNmrTvarJmgESGORuYYmqbJ9Kunym+Bx
hAyWSH7boXDESKWfUby33hJIT8rVndvr0Qc5cPa9y8xXZRtShxNy4gz0qOmUCo5R/CrPxNFQpLrX
t/5E3JkS+bU23ldT8c4nzhF14Z1jTn9ZuIGiJZA308T4XTTIw/hxU2uUuK8marcwihLE2MSnPPeC
klSas/UE4Bt6aqYGeJQzmC7rBoi19LYsA6rXssJ+Ux+N03Cf3xZ+9cjdEdq6kILZZioVqtoVQK7A
UZC/xpHeF1fUjLTvkOdDaUhfZSpIdfwY28dYQdeJsBCnWq9nUCgCbT92HX0lLDOWeUofNOVlLB0w
48w2wgPzBMSvpr3qKXdDWQOaAVmYWTs27ZQDCVexqFONRqpg8MHiIKArkY4qWOQ5MZzNvuv5ex7D
iY44X2NlEwaGaqwduLy6QCBE9rJ8o0oDTo8gQMW+NgbL6h5nNrJZJ0hNZCeYg4BXveWb48fYVdmo
OHqTG18KFDFuJYxas802FwDaFcf9Dlx/FJF3RIwbq1C4uBSWBotb9x/J0hCys1sc2qmxljlNI6/5
jWGRoLd02kE6uXTy2axX3vN7JpSgwjEi5RtY/c0P77XxHWcLBu4GU8Qm92Xv0RuINrGiIPZt0b8K
XLH4krVGySg4n5kpOrIZW4mJLghlJcdbWBW8tXeBdt7uXHEFvPUMlDRPBLL/Xj6ELzd8NLIn1iDT
MQeBb5xbt7CpGLdt6vnBx1vKM6f1250K08WEFapBQDT0cyXCOTYZvjUXHfA7ccI4HwXwIKDHkMrW
XpfGtCuDBa1pentNEszPWUFAQR/1+L5Q5rYJKyjwrkL0o2mr8KpRgZAbMZ75BpuUfyq4s+XmlymA
YR+PJ9JrnX5eYiaJRWe0R5JsuntphJu/6M77vWS4iDEptj5oearT/tOHtjxKkUIqKYDUcCsRIkEp
23dpR4D6fJ7QC9FOcNCqZ5mdGIElRc46d0vakKXaHjyH4a330+LyNjPf7Z8Lc6ecrV86lgN34dAI
sDt8H1UylFujTjkeMgiz5pGEesay2tlEOpzaKtiyUnkHVVCovg5pDIkY1DHrHAtCV6vNei2IT4FG
9Kv2Y/CMfSfKN/IUglHJes/E1Z8XT2Ue8GW+N2zbggMWvCk4ZNO6eZQq/CDml4SIqYnKeybPPh4U
+ERVHrCF8WmXPMvWlQHW7WC2ZuC32eIk78ezCPbcw+BMbGM01jCYW1czjxibctebpkX7152tnU65
JMEsZA+1xhtZGe6AU4/U1FsTlJGHKj+13FEqUKRrnIL2+YkJnDSxt+pg5eDlQZgOIKJTbc1+8iHP
nyKc5/l4/sAbCeyp9P6DXICw1o78sPcKRb/iPq4JmC5jB+iqydZNht6J4UnxcDe3BresgdbZvC/c
KMMQ02nyz7kK2c0jdZtTnGJM2xAB+IKa+JNLMGUemiYayHyx6u2MFDX3MyazrWtqlsom+S4r/mPn
Y2+4GFj6JyxGdO5NubU4PwXb3wOPkDyDsll7l2TurX2oibuW4U2GRoWYKHUFgjMsd0UF1/3fZDLj
0mJtjHue3u+sn2b5I73EVA4z7UHbfR7CyzH2GWCryVVLnani09RrNnUD82CKUl6lSDtQVz0f/ODb
ZujNkAAVGfNEjAI52I/05cIg5sYGK8y/9P+fu2rMtawy07XTfRn3AyIE+WNoGQVoAE1g41ug8KNk
KG7SE9Ef4yeTrifmpX896cGk2JUhrfjzDAurtHmfPcUKV6E/C8hHll3UksmlD3tczSYsqqXV23+V
nrt8q7JAGgiVr4cn8cakokh7AUES9IUjUnIUxg39Q6LlD0fqIXTjWDBEDrEKNJ+Hfht04sSfq70e
J7jh2xLkaxtS1Fzpi03VjthkKoPwq+g8Ttsq5CRYvvSaZ0g+unih2cQvnAIErYx0t2uSqXQmCI56
75GdY7jILqD/ErycOZZSuvtpuxTvs4J1oZZPfkNYKbwasQ6KMfJmmAtJQMvVOZuAh0gEmdELTabM
X5HYa+OX0BCrlYDRY9VKfAd+SZPW5TtJzDaL88BAcWOyKH3Zls/aXjpw195+HgjPUGQLmH9Q2Nm5
9Jfx9mTR+kLnAjWeV3LBu0vPHsNch+zR2sjKMLeDa7QWubGXryJSutt0350rbz2DsBg0Tui4vcG7
ltylZPIax+47GCOcCRTPhhyozvkwH7uHmiGNpiKKA6RQ1eeVxAHDT8adPr5j0fpWEFEdFy9W/CRd
Z7HqfVrE0+1TyJFWQeFdF0lE+AlUrijMrTNVoiCNL0r8YsfTgbUKB3Cym722fdy4oFIO9wM6LvQt
3klH0BpzuUBHfZjy1jlftN5t3dhxs3+O1ci6AkMtj7DVsCPeZ+nr9diNtZOSXmBFwAdVE6dnv6Oi
Be0FsS+zLxoP1m9LMNT7heYxhScTDUqF/whRW01I5pn9PABU7uQE9VUPGLQKzvLK1IMZ88P+gwZt
0ab3HmwtlC650IeJ1Ck2HLh2/Z0GMdciObyeV+GAbtwE1GtLvUmJGnfZtLFWDtD0/F5CoEvleOtR
LidGBKUNHZq52dV/kgQ0B+6Bp41mYv3Zzw/POAv5NDqCgMrl4LZxoY52gXNiu6AAXRX0ULFJ2C0y
IqqM7vqxELOdIxMtpwg6l9kpMpZEYAeWnwjIHGAqqAXjmNFFAKoHJZdLL1zGgocp9PE2yBjwqTeO
ZpCzs3LYimxwstT2azzPBAOaJCfYaHVQvo2tfM9uyf2s9GZGkWswOkeENxCq5XXtb69o4HR1MoXk
rf5S13S3ID+An/noIRSOU6rPBUuH54a1nLh0aD9/K4XekiEc/YtsJXGXGs+sAVmbhLYzBqO694M4
GfvszSSaQKzFKBflhYmhLnC5ot/qmIpkPUQhMGKTot/mIOwmtmD8i1JqLQcH86DBFNqyK+qHf9su
tLdfd6BrSO0S1t9nJq1k+3MIU8cr8B/TwjkfEBhebFcT3Y37b3YDN3jzxWqSC9UNGQiSCSlynpk4
kzuaF4ZZZV5hHX9E2i/z70NS9OFxSVyndJyxJq9E7Nb/HL+7OL1NT2ZW1iigb9zSxx+GGmh/XzEV
38CDdwDN2hFNqn4eDPl9v6PUNEAtx/pDjFI02I//zL2pOoWX7Y8Tfk8cnq0Lk2a0nJl/9n9rqi6M
6iTGZakHbLdwc8zHtnFn4zk2ps54e0eb20fs764nmeJHg6EaJ0juPtj52+nHli7juzynsv8UiibZ
wu4+gaOIFP0FBKNJs2dylfRiDOg6Rfi2mIsvhmP0gBoYofeXEkqCEZtETT6MQ/6xLdru+0rxLETq
ZS2rVLhY204A8/dPWqZLnfD4i4nPtV+sieM6Gw/rc6pwtImyLyq8dMsSm3U6+gdmh0cXzBr2NaiS
2mAXjyzSgT7MUDqm0HaUgHHE0wzGB9aDsIgclOdGyN+C7S+qaVa0kvjCTasyO15UH4nmCQBnzq8O
zum8sIqePv0jIAiQ6Hi86jGiGRW0/JvzH0NQSAbNlqhOiMmlJPxOHCac+JH14Wncp7od62GOhNuK
ukDAxCW1zifC6VGwzxUzh6W9A5w4+wrWImVS/9TaEDhJi32ItLWwoSUpRi4ZSbA/0dUdudOcbX84
t5bzbA6v2B+y6ChVi3PAlcfHMz/JODk04AD5FycZHQcQQFk/f5W5frcaIzjuDsfcT1MjKaLain3S
IZj2DbTlKy9xBXoZttWiCXG5LjvFTAdB/RC/mHXvN+3AdgzE+IcONWhdSb99jXg1HllB2GkZH/0K
cN8RrRqw/7WfTgrw25sQjoz497QsZHb+H2a+8Ym6yH1Su6F1NvSJAhMPbupAx19gpGEFfiadX1CY
aKWPxTAp/EuXv/ezWlnrYSFAXybJHe2oDbxvdpLP/R7ldFMi1GRz5TUNIIrLUkRPw2SOuUw05EX1
DRF8bRuwZpqr96Le0r1tgNAwvCDaEhH1uUmYxlH7qFW4deb+zTd4tBLD4z1OOIrEKzLFfoPIp2ip
OTVEV/QCmphfWa4w0W84Vs86Zs80G2ks81Ggmn77V0rmwegdngRTWK6gfeJGGG3c2PaHowX122ns
iL0aAepfYTiINljmovupOvYQk29ItQwmxgUKaX91LyLT7INUjLZ3gEwTJdUhfH1DF6gtER6SbkqD
LgDNPFTYXgUjKY3dnUPaMmHvpXipqfAXlKv+2klNIt9mvYfm3R4aotl3RBn0J/eW+KYJ0rRQWrrZ
TE6OftMzxzvhUey2rFMp34BqXaJHQlitamiR81dXdDiLf6t82kOlp3uh32JsLsOuRjJG1P7HB7A2
A9On591ymctAJPb4lvU4R91Dma8UZ17ZyBDqeY/UhQTs7s24BMwWJsJ/jAWPc9+eBj4xOleBJAus
CMCXGVcWoyr5omRF+9ZlvLMSxNx7vZnNf+kCYsqB3jwM/BE3r7WIOAeo1raGDUBApXj0Aezq7jwE
Q0a4im86clOeiXfAg7HIrqbZCL5D6j9IzLZ4bxNWgkr7RCh5u3eJnkvmODBavVSt2WVPHoPY+asA
zMJKndLCygXnJPFp76C8ItK9gGqbxaifA0FG5hY0ZwdXt85c7ZVNLpWSRNUpsWqzIGKiicWMU5lF
d9e9s5LM/LnaIRSceD0Jyn+mvhxRPiQUXjSD6ipCYf/V2pOeV6r3WhPAOJYHYWw4/UAUzKwo59tC
NTf6J+E1UY52+UXPEKg4QDUQym23nveoEsJM8rvYwO2k9zTb4lxdUMt2UJc7s/Qb/TucL8HyL3mB
641gAbm4hLhI714QgS0GsNJKOIJEACFpkWW+l0FdinuzB8DfBA3jvm8XGz0jOZHWiTkX0/Wx6mb/
BxC26EtIFKXJFqFl7SwR8QkPCtARnnc96+DJ+wkt+kXK+WekSNdMWeyJntfTfzyf+BiCmnekCPPC
bRVKhNMgKhwb0OezzEb+s8hxUrVsg1YfUiTo6EII3n+i7YMUrqHoB1F37XY/Ot8jQumGo9mhriM7
dfUD2j0y63e3Rg+ZnLGo3aef5LpetwI759PrnXZTMJD0XjxgduWE58RgQuOcbNh6PceL8yaBYaCa
K6tybxXjk2nOHnXclaY3FcAry59Jm8035upz7V981pSxUw9z94VymZiLRB82PxXnaI91cu+2GsF/
6546pU24tGwxMkTwxPa32F3nrBKglLKCRtm7m/Jz6q5Lflfz7lMC5McmCPdwuoms7D69N0u3LmAw
RcYCfFr7QLlFav2SG+2hjbYAc66B0WXrvMALoBL++k4BGoufLFirjbCXc77GPlMyrlkRnpLRQCCX
DZYL19UahQgBCbmY5Znh81Gz5N2zi8Z9KvIGIZHj0Eehu+UGbDMjzKUMkeJHvI9JEXutWTwzRhTi
ghOBhVqjfi9WbNT5vnZMdip4fRYJqYBsx1PvpnTb+TH/DllsSCHhb+c4h5Y3PR0S/Fbk0x1Ayd6N
wP0ExYGT3EMccYrJx+3PTszXfjmq/MzJ8GbiU1tt+7dLBm+jfWAgSfVYvJHlUPcgVu5TWlaBW8th
mIOJJfrClIuC1nN6ldZdqn8cHhoI6W2oj7ggoc4UAWbRYt+l1PhzLgZ6vSMDpeeWk52PZfYfqpHq
y3WIlxDmnU53fboSBGhbC6L8v5uuEvx7ruW9WNwY8ED4ceA0rImUVIvLua2wS81T5TvX97mfmu6n
Tlxj7ZwzK8mM8gnFJeSH+2SluYRfhWmdnHQ2hMnySOwI8dZd9rslbHPpBR4jZs/fRpuLOI9JgNmB
84BUFMETWLfKUhFv6AZwqqptBEPp5vINtfb2uGOnf268MSN/o5MLedQlWsieAiSTKHSTLr7Y/xEP
4aykQTEQnQQqrgucp6CmyLSNTX9tbti1Qdtoo+oqWLt8zTsFN/lrm/tfaTeKlseWVkgSFzpLrohH
xLlj8JY2gZ42W5iUHKfH4XOz81eSrEic8odXP/QIE/7bHipz5S/+0A1ughGo/PWwH08PtN1jgcUg
LslKhlsX+yIBa4dr3lY5R6oKa2cNxgYMOxEAdPgKVLBdeI+ePy0rvGO2Nly1IfrZuYDkThfsxmdE
92rMUnWkrofYQx09ailmg+suWFd15J440i3eQBPW8Pc785Y7WsKQ53a/3cEZDunTftdEzFbS8R2d
ruuDXfPt9LJyO+oQK5l+T+oIAUqm8wjY/PhQrSWIq2/uqdUWNxgGVSCMFW0BvcyBO2crYg24Lmtd
ZupC7og6KIZI3yXzS9vP7LuMlGsOk+ewnLwXeeFGzkm4iqqICMrm+9jCRtnv+t5K+o3y26WyOrOX
w8kS+DI9WJAvo9rWe80GN7fttbsnNwIi7KWDYMUzKL4R25+em8+qQNYcoW645wFosu6pM+X3GPiq
Tirhp9HoCSEv9JtEgwg87K4NPcA5B6t6e66ScOypJMlWdAVvnhOJFzvyaG3Hv/3ssqqWxqkGTuw+
mVb+8HunSO8BYdfuuLvQUjfjII+okh1eKnkPz2sG4kWfJ5LMn2OFZJ+Gy43nHRgnJoT1b55eUanw
/HuKPV+omlY3SVhZA6Wwz974OgPQ/npVhQBD9F17d0LKfBqpXUEquwOl1J46Bfc1ekH0/YphffeC
bdFk4wmuZl0t47222t81wCJezB06KVS8YM863wxlEeanQgUx6i2tkQJR3aPFrnF99OxDDuXx/VJ+
Yo3f4wEVfSHeAwY5sgAzfL+5aIA1fJSuChvMaPCxrMtqN4PsO+QYJ3NaGX5wWsQUwpcFiLunql6g
MUI5mVcGf4rxd7L/9+E7+hAeaWagAlGGAUcJ2EcnsGt0XTxZzMEChllFDpSxVJYLSlXBQuZ5Mwsv
QCNreUn9hpqcA21HC8l4YAm4OhRHK6VEMYbspMf9lKhdjf7Th3fVUJebT+gJ5U/UzaabTyvApqW1
5Ob0yGsOZHngHCRgPohv+3hFHGlGjCXrFxu6UKjoqgW2J9R7iTCjbNDVaC1OfWICGeqq2jo9XEku
XHch1ZnJppvoAiiDcWHN/R+2hUJCLToCD9/XvXqyZ19H5Adlsc/TeOvOsaudQ6q97Kcj+qDu7OWz
kJT2baPSzv4iayN2xXaKNrMDLUOIp7Ax0ulw28wA4br1gu+DOSpT1JK+u0Qsdley9cc5N8/7GeA+
xDU3pGcRVLYKhgjsrKpiVXTuWja0sHS8Tb/4ARyq4kpuYj/eNPcPOj85olOXMwOvoM8SAAck9hIh
DxmuHkAPaEGl4hZwTlT6+X26ugGaklu6IrnXoS/ej1nwXMd+AFE89u2VqFJMGFI3XWpIg5kKlb/x
yIJ72NaVSlEeAmChvfKc5LJtw9ILewsxJ7QCfNYThcVLPRS1qfvaCyHox6s0x9adAoZDDLMmH5Rj
drzp0CQQSg/Olx38SsW329ZGJwaycg5OWhX87uypfE5R5ZT8I5GsLkGmBBzPNOSfbTqgrTnqylRZ
mxYZYe+79YwPZa99BU5Tf2845TuqaCRRwq9vGZb6aNt597bjL8tdHhV4z+da2yb1eNDbvenLQoSp
nEejGvbWLpJoUXgGGnlov1smX+og5ZXzQYWw2hR3kWzhOVckruLpEfyxo0vU/Y1XKwMzCAa8hOxQ
iwp14hoD9vPBS4Zwv2ldJJHaUpQXnS+Xl6+K3FuX9pDfRyNlz9ImklnLsXtm0Qs7ZMS0u1r88SBc
0NR6t4gk8EPhdoiLk2GCKyYnPlOktoklkJfxwp7/DDH+ljnQ603X2B7vgwCdvv9bX+1hca8KKlqZ
GrAa0PUs7fvsApYhszM8kcrJ4DxB2nrNeF18huOyTLUtlSn2h9MjOZ87OOxY1EtN5y5FY2SCYaGD
o8Ppgk5Qbtpvhes/DxjzyVIxoD24qEH5A1KgRI4Be/ldWT7LR4e6nzdmTB+gv82jzeXMa4t4jr2Y
uN87mxYvYysrqYAcCtYcMWv8EuermgBLayuvLI8993GL+oJem4dUieBIltCKFZH1NT+VIU54dEzs
KrZlCQPMJPjI5fIvtT4yyJkY4wQTB7M/fPCyqW9EHhNotEWZh/94z1mTFkTx1bH7P+6IWkemQApE
c6DeW98dtXXyXSy20aCH0/Rg3esWh5Kir0UE1TFy8JBndu6BuQRiEhH+JATuFT0ifdfh3jlPLtkH
3E3zaqVNnHKG39d4s88dcCA+t/0iGOX8mTusbwbPG+04PPDmbC6ZURDpos9B9I4GJU/nhuoKhXNU
kw+OXbQAe8NGmGWlIEsKhmMydTps4q8EzJHWVOUSdBbBJwQiWlCd3g6qlZVUn7l4D2i1dCXsndER
zTYOA+waROnb7jyXIYqOagz7DIKwMmG9VqWvkVmzPBBmOuwgfAS2dsTOK0YOfwcrNeb75PPMa5ng
CVqKHPVegIXkXm8YRyr8u2/faxTS/if/xvs9XamkELpdG13m6zrp9526MXuQk/jBPr27+R37nGmb
uD6dmiEVB4a+8QIDkeGxduQrcumTNT19MxZZKlZbyMw4Ss9FQCf7W2BF1EterzVEBX0hl3PEvtBr
SqwDPCcH3pFs2MZb2ZsnPL1HmCVGctdy5CjvTedte5pCtOJiqYnV2ED8nRTTeRIXJMb/hRUrDdLH
qvbzWMXrUXPLYVA2IHvXyA4/OQGZ09/trto0E+V720GSAhm4rfhGT/TAxGRLv5K0jUgfo+f3iTr5
s3OWwLoaSSLkCbveyd8DMSuiBylCrByTeGfgG0I515rWnrNfADf9pTro+ndjpXkRYAgKBQwOiZy4
etZzC+UsBUTqfrz9UY3CwxA4sFkZXjAbzYGtwbxb+UDIZsHW+1L5LmlO1WW9Inu/o9O3rFuf9w8x
JURmGrU2cANBtXOJcRWuJY8Vy4o5OIS4430ajQsAhXl0jjbWYEYeKoxsRM+p22qonEr4gOFz5TR3
7XXoob/W2cjIESTrlMZGtVGnh8mJRQ44s4Ck6NMiVCWCATzPeVr+BXYp1QSGIee2bkW8b02Yop0P
wwzS7wdgMRHrNl9ZvLautnA903M3dwLcVvRrMuVdvGHmDI1/zrv6q/UYc8rBexSr7O5eKhtEpwYk
XkRXFF14PUE1ihBF0dExcyiIkHFaPWBYvvXMxGbJKDF/E8QsW9gOFI1qjQnZj3QVzeN3OB8+JzyS
1PWVeC62iT7j3a1XHkBNVagxUzSfMehJA6ew/xBFPbB0jlP5UUcBxHaCtNo8N3i4JnXjhH3RX0Ps
pT5QtWgrjDGZVh0ADqBpNHS/K22mvG+R6tubbF1ahFTFjV68J8muqDNTsQfM9vUP0Z0vuz0UvyI3
J6GDfnkANd7i4xZwMj4tWetvqliMNe1N9oyjQfeRaYQWQxAqSdjaI5T6TNyH47rU3p+wONEw6DFB
HsK77jcJFanAjxqPV4C4Q2abqjJKNEB/O585Ac/V9Vv6SsOVR6jykcvGNkMICPSwUuO1CxbfwrIZ
+DehCkuMXhSmcr9QFQUd3rurRRZ8FBgeq4VA/Y/b/sMnMZPauKGlkIPbvYwrE8zrvIVyeLSisII8
1VMkSqEO4kYe6YSvN8p6EzZxfEmsKljqNxMPiaTgSzGr420eqrmuSE2ThT5G18gQEteaTN6fgspk
vNguQuXqKmoRnzu5zCrZWxJJsIZ6jYWmLBJv+WcLZ5OYSQHsbipxFG2ePSIsR4a+0mjruPsowa1P
GJssTdqTvxUVK1iVpjL7bH5ll3G/XQvJKbm/eMKMGn1FhZN2qPVgyTIyc5TqoGHs5m+8asMjPbm+
g5IaDZ3U06zeAIjHPztvC18Wc14FwrMlCPEMeGfuXyf7LN/z4ltY6I7E8kTe1tV9/lgFjtmljxiz
mjyYVtS10TQNDxaiVHwCqRiawDzHUr+aId3h7yk9k29Nx2jvRyrdJ4Hwq2szdzQj8hpxV7YhdFNf
Xc+YJmMTzubEA/pp+t41Ik5juGCp8UQnLbXSr+laey4Ss3LNK+bTbJiEroUcVvlKRhv7grUe1/ws
QGDV8gQ0pQqqd/Ms7NMfdNcJUP3M67nIrNv8tKasp3k2N3HOHBOB/u1T5dy7U3yovknAvhJJkPPj
6a/no1Cf7RNmx6Ai2B4uNVikrs+1ZY5c2Jp60GhTpvwvYJlpq0V+nA8jHXaOhgavRjIDD3F5IYQn
bfoo0npV0ErlR+fH/hBfX9zxZZh5ePXCuTHsfpuWfuZJ49mdfNI1JU+0ucGPxEf7WlHk+Drt21bp
rWApdaWADTiARAP+5b6VgaMvlbe2DbtMmDuem0yQ/tchjsFcx5vIoTvmE5MMoUV13N10T8NwkVGS
y36hlq/gKGNuaItZLGc9svdhConZ3z5wvOQXq+31KhemGhaSIwJV83nh63J7wBncXDXfPjYRedDh
VZ2aHvXMgUQOoEZe+RptuBcyeI0sDeQyvqkZc8JcNaqnb7T688qB38eIn3v9fWUB0gQfv/qrBj0E
9oZrVyaoRTSG8Qm/g4w3sS/+rD4aQwpRSPjTdBnA7f4Uf29yWbzHq7fTdiaICT7pCkMmUNCKRmCN
WkC1I9P8W4OzYp9L1LdjO8ybdb68P/EkVz2Ku6mYIZ7GDa2yFTuQmXXY1RYMOSSl/JE0xrLD/+e7
2mq7ngtLzP3mclSY640VMMNS7nMY0ib3iyPFnyt/IvEhPk0wofe1iYcXPx3gpqU+BUYF9qXjpYCK
GZjebHOg8fws1erugJWYN5CJNK+RJb1m3z0A7G9MS3zvYIYWDcGWuH8shmqReZMAX0TI8haazvlj
pWZzV32zBopiyEwSrmA7TzDO1cYJDiKAK4COqElf5I2Haabq3iIiQfSr+L1EnwEif4r4dRDjPQec
J3b5NEU/TQavFfjvpBDDqNGwjlSvuqcXTmkmBdPNuvy/xtg1vNNDgP/vxapcdSHGHat8/xRHknJU
ZcZi5yGzI4HFicQDWcc2NtxJDCK0obHi0R1BDuV3gE6O8l1FCsMoj+sIb920Yyvp0P+/zl1s4yeA
Jc69kC4F/ln2ZcaKuyipILaZXgTNoxGeNqyHYi/8PTwoHCaBxNUIZcDzrg8xoLize/g11xmxyce+
6ZrugJflMjajyKXPWJep+dEOoe+88BI7AHnh+Xec+XzT+TUbOzCtWKQ8Wrvm7pmBVNU9e2ZMaDVC
/42DzvkoMJvpEv6txSj9Gn/Jo5or3NVHh/mfPhDoCPzqTEVhMcj7SAIfU6JByFGGLLbB3FsJwmsX
ffubjBaI4gfLq9a5ArNqH2eog/I4kgfiVPKVPdG6+PyJ2VoXcfskbVHxM2zyFLTzDoVk3xekJYF+
R9jS279wE/BpIs79qxISslALjqgNWbHnZtv/lt5q/ikamuYmXvOc/zMTTnM8LRBsiO8MmgCk8422
W+4mGqY5mQOJBLxfUeC+b8ZzEKnOXvE4Oyn7tG1qr26HhkWJyVpKfk3bNqpTceiiYbAq50mUYpa/
B3G0EFLNaC3HGSFuPs0Ije7ghe+pZxKZ4gf1pO6JfM0cNy1fjTKQi9GUwc3iv7x3ToQbUbe7IYgI
5Hih5WwyeBI+QtE3g8gO/pbYN3Wjiod2mzAl1ROGJyHq9/sbj6lyBmvDUdDOiDBK6eMadDZRLDKJ
ChaOGdE3RKG7RtgFUpIrLcIR/LDDaaz3Qx5E/N3jNEkXYbCJN+MrbA6/Qm2FrqFRx3ftrJNtbYUe
c79TOQAsMx0R3o3taptYt4thcZMjcj8wEwurgJUdt/OOSy+qCCuhwDK40SR/MzqsWnZyfm+I9IoL
vmysDfREieW1qDqXIE21SGFgJ6SHSHEj0zen1OQwX28fms6LWEat5X+QLMlcDGrtrHn+DRWA1QZF
7fsqmhCBDdKpHLzp4MtRtqmEC0C+4Bmp3LrVXUGVh70KqZtiLv/kH6hkYqv9SM2VmuyQlUmQsNAG
Lu/4O69a5WQZXnDOeQ0VPYk9TmwfsqaUXOWdgUzXbxrOp6cqTOBfVf6nTXnrpn0VzGryxpPT5ovp
GpuJlHlri/fuKxv5XiQevl7X0ipct112/dlr36pzhRl6C212fvZiMEUtLX1xqHp16gecFBidrJzh
bHxnG71uePiRmnOn2RB5Jw66Fpsvu3/UaAkGEKFC7VTwsfBwpshc5pDdPiNnSMswkTpz/nrbrfOt
vvMYzag/kdBtarf2Ku9d8A+z+LZPXOgsALNX6BWusqdIrlYXxUw+61yyAyB0YcWarTHjiyHGV2dP
8WvTHkaSxN5YM7XYabWQoLX0nCr0KQ3I3Dh0FZ4JlcNKqUGnb936oYsVFCTjm4yZXMQGl2PpnlWi
1eDzuKKUHzvL5D7cTKMGqomFReJuJ/GnjCwi4yJXP2UhAFWpy9idSpjeGjAf3NE71PizdvXb7hLL
P2Gte7CGolJynqV5+6cb+PBMGM2WuP5H1Krf9wBOL2Q1zncznDxnVLApZ/bjWxyaZ8qTvK7elOJN
ym0xhdirhm4F5UMSpZbk//7c7pI6Jx/oUH5YPcJ6DfTgAMr6bZtLTazTkZs8ngDIDRnz9WXzqQd9
TMgd1DoDnb2YIUh85brvaXXfLka11foTAp1891akTrNmfhEcuPTzyXGRNY/NfO4TINMou60DoiNy
d34if+Hf53Fxj1qpZpd/chpmrBr9ED+xnZh8ZV1Q937K3A3mCqjypYbevsUDqNTu+edbceWjsyLA
wFApRqjzsfVap4E+y10D+HeTnl5UY9Ts7cy6H4EYr06mtnqfwLrdCLIARWbOef38aTNsIEmp3bdM
jxZ3zVsY93cF/ezg72k98jowv0qJNmDVIet1AIrjsufH7wnHqCU6zrKfHgRKrSM55K9rkNgo2nKG
ifRMYs9ibyDqvUZCVCPn9wbb+2Xnsu5dtFQmuikQLeg0upzeMUqCNneywsdCdlxoennJkHXnqnQI
UcvmQn+LbnfbXuROeDu2cGpab/SSO0pjSuM7TbZgNr+cDhF7NZtfUFoO5DfkwVSOlwGNdUxhEFLY
YcSKEmtfejFFcPUVXiouZz6gcOJzYVxguTinTzRxfzLs3KiUIAissuH3KeWK++fLifMdnmtqSWu7
r8slUc4OkNpAn92yOLBxbbiC0AGDSK/FZ5ysU/rDSBviCobMVb/wF0k651VQ0qR/T4cmgCjh0kTa
r2xVNo7XUMxhMpr/WKjGQ45pNlquqKzeBq3O8MWQTWHYpvYK7R7/Tyqf8DRQ7bEn2IoV3Bqy0bHN
MO5PUa/VZ7j6neNVfwn9VMqjL0IOda24FeArQZRSJZaWDmRGZ84Q8QbeVuRHrsvq7wcNLciuexTt
YNYoRzd7OdtxvjLbRhlkD4a4IwLrkuTk29pdaX+pzUAFjN2PO7jvMXw+u1Im9DTLsdLOXTfCeooD
vG56aADXeehf7qCXO81XHY9Q+3+VLSef5ta7bJbT2QW9uJ82HYDce9m8zytKn14lOQC8pBJSxPF6
Dfo3N2CavMQnxU3zUJdjJjIow9cAZANTR0XzhjAemQQuAODUfL69ylYGzhXKGfQquqpFRp0BtZ4E
fV1foP6POTfiF8pgg21bnhDttl0o8G+e0QrlfzLLGt/Ed2kanVfD2F189fQsF9ytxcIv2gfkg+Tc
XllCoUl7C8BRJsyg+7NBda03m14UdVuDRFKzqBlnmRmJjXZT957xsMEHPv6iL0tw4y9jYOgsDsyQ
eFDPWJnE14oQZ+DhPx9EoxBixL7h+b+9gIJjiM7OQQFx2obj3K8PB48oXcT93Pd0VqfX2JxT7Ar7
7rS9WBpFJNKgfFMS3jpIexA9mAGo1mIhRsRjziasMYE15pKkr3yyT3bZu/I/OW2nJt10KG1W6jvS
ecXmr3419kjPItlDF2cTZ82HQddzkEP+XveMsuYvxlRTQ9chkIltZPt7rMrWNRwoExOwW5noZgqr
HtCJEV/BdyaajZ/CNYO0iKm1j3gx6TfuWDMQq56ZvC/7uPMxPTwsWCxucbhOqdBCh17KFontOH+8
Y/E4O2ktoVPLB5QQMO17twX9s2GvDntAq7gGp/a7+qsjVim0ymbza6euUfTj/n5MpY7+wBouiFAu
Yp3ZRTrxxx/vVxDW+3vrd0DA4BTtr7NfvORU2qUjl3SdEG8yYi12Iwob4SOnu7JhN//6QeXItS9j
0pjLCxDjKUOuaf//QhnShhGqukMpyq1kpraniHMhjhE4HtTR7V9pZq8giENvAphlNIfI1XHQ3GSI
A3JDOzwnTKvUEU21m81Omh1lX876VJdbGWJ6cXSq1o35HJKMkvMIcvc0RNI1RvEUOBkTAS0CI0zc
YE6NCN7oTsYO20rK2lqR9XmLxAiiEZ7C9TBX8HBOkHex/EBMVB8btRnpHtpxj+ElIHnzqZGgMx2s
vAQdJiNXS+2cwKZUeNmmeAP6VajUz6eve3o6TRCtfZTPu0dqIsMiTTOa5PeAxGRSvk28COoAn8kO
59OQfYrfxRdFkSrtcJmn8WYWlZ5FaMI98bTlYRv3cFCVr4t7ANj8JFGTmxGppXf78Eg/8e+KnIRS
cQL4oQ2ZPqF6r0o6P6CF78OX4RjF0ht68Xepa4gAaHO5RkYo4jsTe7kHR6YQInq3jDJjL6pMUkOo
BMXo1GO5G4ac8HKH7M/bz+GSKx4Ktgkxx3MVErgeMWXk/Q2E4U8PfGCAKi4KKO7St9ZGNsmGdLFd
O2Xuwf/KlF41+h/srPGKUVYdsisZb7Y2gvrZvbTOLQeMY07AemIcZ7FqIaI2/Uqwsm/wYleYK1Vu
WgHVXp8+99gaPydfEawC4yznWiZXhjcpUbj37kfatBNT4JVp8iagQ8zbJ2SI97jhwxeVrU9t2zoe
ZJm7omnoPqaxnKEzlSH93VGVcTw5Mods20MNjY6gKYjlhaRKB4cbB2BwqMdtXeLJ87FET5/Y7orT
fSb1aJaWakuGR9zo3clidEsjc0H851dpe1KHGobcMzX8uNS28m0IFbmWe+7JdZjhv7+dT+yMTjCO
x/TNNDt9M90rdtDiZkp8AMhquX05L96sJ6/QzRiI5HVKhFjZA4h1XbVKBhvxo2U9vk0CWy7QODAN
9UC9W9wKSpJXp9CWi82aCOGtCV6azEec87QpM6FbCLQO4NKx4IKNN3WsQFPJYlrBjnkVfA/9oUZw
3LFAL63qc3PCNXv7Ipa3/kdRNLsjLIkV5s9TyNcgwoxDDAdYIkDUXDztJVcV/6gChyAb2yWIluic
XNMoxSP58/UH+/d5Nd56Rhd5m6WCNbkIKyeK5qjHSRNulDW+hFzxk23mApcQQ7TiEbCvZAgQA45e
N3iNuhGtgcBhEByTfKnNCWnbmUC1stjghiEy4ncB0ViKExj8JdA0+5GuEXq8agR8JCgFO1S8CHtD
GAhOfT84wzLs3J7QIhJa5UhsLPNf7Vd5aTKhW5gj3a+jDtDmVaJl9CWG657q/GPyN0LKZUdJrhLA
bBag0HxFe7IOFSawG/tcdR4rcnkRgIlZKHyQml1+NfGk/iSFs18tP+cBFzwMz9QvLycU4HXj5Zz7
JkEERSs+ZRjCVeV0BbV+EAanx1zygUlrbF4V8lrMbIWkUBLvHix54H2LQls3Qk88uwkIniUn6M/A
M31Mzod5SnMl4orI8ePnWOUBAZtQcZyf2UJisw6vRnKvOV4/fxcjJUIytcV6uW01cS7R97jnl9aN
kuxpO/EXqC0hUk9Q3ZmjTRlkMXxxUlNT6lG60yvKUjEszT7P7IkiVGQmoc0nLje51o0SSjd7nftc
F0zNOarz160DRno74pnqwoIJDogYzocttkZs9hZNpY96Xds35Aw8EA8gSjbifkt40Zi025gCfwp8
pQiENU47meFkDdxXk1+CkzlU+SbV0RvV3FQKllfdf7M0ttoeOVops59JjJkxWN55hdnIx2F9YbSB
NqIvsE6zieQr6gKGpdoHWNesniqK7i5UCj13UyOODMl2r92IgNJimdTuobbDnE6HgPWWrrHhqW1A
JUI33UyE1NXN3+YSRlrYVbckbZ00Ic1GIHVZuQS2Z70fwz+gAmLO8NqddocTd1ZV9wldiafrT8/a
eYZPtokic5fKm87jaOFPZ3Jl9J0Vx80IbY1kLkMf/7H95v+aLSTLNfUv6xBf0LcbLcKGp03QnKQP
e8/P8r0Ldm3GAhH7M+W70qe+ZoxXrFnJ1POtBwSqxYeLI7dVSHQVwQsvBEM98Op1n40qrINf/Vd0
8VxpXyq+kORrUPu1n+zcs7z1KJv0gSvOvPBIUU+cMBtIuQ1cDZvf76OWwko7D+uXxQs6QV3KVc7h
ehgEUO6oktnCnnonDZYUfD+ZvOXnDPXr/9KEdAm9K3hgGFHiKlg86fvirIQZFGp8bFZ6pRohMBV3
rntJt+ZBAFnuzekl864mNZ3E2VocYF6rDqV7za8W1VmAYenqczikD/ow1KkmzenTxYZn/FK7WulS
bDyu6cWsdr8yiDDy/p/v9fDizDlzcVhmLeS22/XeFHPWat64G3IuUL5JHv0DVo8J5aThZtPA5MWi
IPi5GVUEEtXMrziNlwM+tKacdL/5xI3JWbrHfd0cbLDCFZXeJVPYaxFYxKHFYhEvCRzXpDqCYNXz
ZCOi2Jto4b18MheV04NVhiQ+uDfid3QQ/k13JOzNuyxPD7Yy/IchIIYN46XF5CE2/komASXoGBQG
sHn/foB+yIzTlxEUBBJZmz/WNweJpfKKkFPqwXeHXpMdQ7mAhnzzczZz1KsxFPJw0o8dj+XcPIZb
WgxuQYhjr8x9iwCJ+lY8iH1YPFb2v3NxbG5eRUWcNbLWIZOyc0srtB5xr4xEaUtO7iK0OlRICf2y
2nSOgCcgM0RMvrMYw6SbdqF4LAKvyl/5d81TSZZMHhKa91AsjRppYeHU1RNGkk+zz2Luo2xdrBea
ktik33xcQbBdpKWcf0VdT4lhiCQDQaeST/qTHh3EfxkJuH+L0Q4y8DVkUWE8QGYa3eWr7rp8MHhC
ZMBXvaDqyCYqNKG1yvUwKoudaLCwLQat9nC28PceSB/CBGCcupXziXIlZ/eQ7mpQn+LgIwIFNOG4
B6/pm6G3AeByQGBEiO09wi6+BYilfM/johP3Z8xXqiJ854aME4Dyud8CBhZ2sIXWvWy6IGCzPIYu
7J59lP3B7ylC1yCv41NdjsqLZ7jd4hxkzvh4hV9juEUeV5xW0QaU89xfuu1PEiq2WIybcylcmXYT
DPSBhnwrmmvxVTv1NX5rghhddTY+XAaW2Sh0vrBVauo7cRcB9m66ElPzD8l9l9BGebhSA0+MTJsO
FvloMNT8ZgwKk0ClpUz0x1NCYbhWMDigLgM5sG5rOIy4XUVDIK3Qh1S0mK35ncz4zNFG3fACPPn5
2efi5QIT1VioEpxUd8EEXDj3ScSXq+hAq6uw3xY/8ND2IAuAb9H0poOymLX5bPyT00rPxSLiKvWa
eOqfKKdqeEnXyk1zYz2Wjzql0R9Zct5mcMs2rrzi8sykgpZiEu7NxTHzHIRv+LBLgmkH/O6RCA+G
qCTWk+ehVVioUyUQdcb+Tb/STYjXcDrIjATLFNFG78if8CCQgTrBkU+77kLhRDL6zVHbPCqNSLpO
htXbmS/kTCx6GbPxCtb9GGmCIXnXObGF5m8bZbSIGf5SnXRPqQmlqOh/DLUAq7oEFl/vIqvoUAcv
J1ZP8aWBD/ypBt75pN90pCnBP2S4brSxbpw4Nmnc6ppyPlQsq1eudbRgSiAWh9pbjpePPP1EVjlx
J5vVK34WvwuH+G9RPndPCGZnUvnlmHY6uoJVv4exfGSBM16B1zoXW7yyr2nKEC+LwZLFY/VMBxAV
gi6ojxt21akYLrNSgA41HM3JRt9pZ5LFsRBoapr9XB0ff46blrwxdtV7iAyNZTUZKNpFbDyM3dgQ
GhTk5FjXgmFbzFjErWgxRY3dzXZm9Zb28yDYdtmab2H0sp7h8/3TQ1CKOHKEjl8W/r6Yh+IuvtuO
lTYcpr6t6oUgWvKwGnuRBg/upjimBGSzidfbhv9urcHBdiXRXsHn8tE9bqGrs++a1BhUFnrnJDpM
uax8C3qODZjZPE6LeDM9jkP/XWTyfIwZ3ruM2jiotMar17p8t1qAWJotL/UGNN6IxlwZntyNTeaN
HnbUB2EIKBW/RpmpoTuk0RfmZ41br65W9XDMG2E8/LVuWCa0qaRmoTtrYq+Z4fp86kqskoRu7vQL
ghwkKCMedupts9d/FLX3K155sEeTf5NIiBLg5PSj4nc9rLcseB8QujtBR8mM/aMj4Lq9cdftxpCv
+aPfN6/sSBwxCZqcIQ3Y+EkYeyanjga7XfdGIb9WxTxagvmP7XCIU2D3ztdcq8xzHVMFHhEr12c8
o11baaQmZU1N/15zKmsNdT1ti88r3d1otphYKNOccG0G4eEFnGT5Nqbv/kbE9ZJXii2dd0vqs07G
LAFd/HW29ziMnScS2gkhYo3XyphzPNGlS+4FgqZYydLF1/UqbJSea2P0JkNTrf+9GDYOMQRsdIj6
Cr469R3l3z2Dtkc98xMvICqwd5RqVK2aWMc024vEmdcbj0CQt2U3BOuKtqpmWvn2AOn17gZQtQ0/
I1CslCogrVGzQh7Tr8pfUa/jKNZgtJqp0rkaIfeLSlWSNyXu0KsjYXBRfslpT4p/WJIfEruzXII9
MNjELhuK99vhLDdn3WHVPltxckBSYfhtF9msFcTR/r6DjQ23jxeqeupLFVAmWVf52MI4515z6Ugd
3CYfOPxD0CSz3FP1bmZ6vUx5NDRm9R4XVsHAb6G1zkksKorOAIHMnuRu7OL06WgyDhVeVWS/Wzvs
FSN0iIWKdNkbYk6UONcQm3f9zlUkHrppLzzOvic1aO5Ri/CkVhr0rjtvC8RpXLY59A5G5AAfbddm
5d5rozvayFZry+12A4QnNUvxB/F9zWDa4GSjCpcjUYOHQMgraJBcndDcxPK6/zhjMGcqhbwSWZ69
rRmjShZNeW9l3PiM+qOC29B8Jrr1QrkbiIa4a45ueAWOCaq1zBtd0mU3m7eRfGfsocCxi4N8OU9l
8y+PonnY08WwBl5+ffKB2dU7+0f8pf5Gpz7eQcbciPMZgK49dzBLmEqxtm+YP2d/ygk+kHuVVMbC
rHuI/e7Cgol9HxglA9ypmkZMYbc0ZONp5utSq/ohlKmIeKWsea92SUKd4RmrzMTzdIneW5FsEzUB
kNFSO93PCoCpkpTT+i7UQPBJZAnqeDup6qPOq2XL5vEcxYU0ISgANwdbst5vnxCYJkwWUQb8xMaY
VQJ6fEKpfLhig/XOLQCOmBbEWYPlUNplh3vGlT9//OAtOPsiwzOldjJDTpaB89SAnmjrdF9Y2YVh
tXyFPccIi6V1pDJs+VGvvliYvkaVorLlG8s6PrMnQu+02YER9odR/PdFtHMcr3/tRnjwIbiYqgHa
/1GIe0bkZzt2JmBShvCdXCUv8YjnS7dnvl2lYzds+1F3RUJLIEjZjBdFG2vwQA0PEAOUGLkxFS7m
5TWPgyciON2EgLeNV0YGkRaCCEjJdEP0AIuiPbSn9blZTgGomjvPtqWRC1jelTiPG1LANqK5eO7W
f3x2TahvrOdj9lS7uuERmF+ksmKx0fwUvL5j9s4NcFaogn+3Aolg0lG0RqdUEEdL2O4aRj5+12wF
7sbCEEfyOjIamFqJcwYcdcgMqCbJrPgrA4QlOqCgheQAod/jUqLVXRYNRbLnDg1OXdxFdOelaEsY
5e9JS80EnUWDZzEf+WwboT++AiC2/sglCqdcZDLFtvySKo+JO7uFK6+PTGALCZ/YyJ2tBvz7prQh
TygLG8ODUKWecF2dMCn+hJEGAlCAdN493DqACmwfYb2goXiEgcs7xEZ8M0JQA154oId0/iQ/jNBJ
rSdqAKkeAejc0YxPykKWSB0O9ykZrkGU40qAB7sU/DtP1+9PUM3IelxLHuwkk4rW2JanBBm0Rkus
yGrWIQ6ylkpNbLXuT11Yc+0DpFyAzNuYRzGJrjvvxfllvlilgZtgKY5FOCiolBuRI1P1rpP7OsYl
GhCpDqLruIQnKLpI3Mk7yqlFy1M6yNxU4c/gPb6M0GXNXe5Kn39TqNFb24LGwlN1z5QNlMBVWNXf
uGnuWsXxIgXG01wyVQ+FKabEFXnJs7rpTBH2wG93i22KLzfaAxG848gzh2zL+s+JTZh4+JQ4gD3N
lF5Rhuxf88D+SPXpSIntPzFplzWi0eclRd1whXDP08gZB+FGIBkfV637Tk/2eXoKxnN4/lAnXrWg
qCRcdEGpMry9ArDCoF9eTobQqSfWBnfgAQuN3SX2XCpOH066DhdgVKAiVwMiK6GYeG+yE1ZQFyyT
8Qqp2j1mkDF/9YHDFvdQxzkQV2nmMn5mh3hD1nsOB9w4lPHfMRaQ2ERy4pbQaw/5gnJ4XEZo9dhu
DRmnrwhPliiMYWV4L6XsdjjO4Ech6u+VosoGHrXVaXAROfeWtXqS+pfQ/5XpKfuYrVQTXYZHRzhn
liQPYo+CJpB/H+yL8sdu95C8kW2CSs2o94ILYvnwKRlZNSXTn42yfK7xVOSs1rm2fxLnV/rWmmK7
B6+YNPnMkpQ/jakSYr8xe5SjTPSvhbwkB9kpgHUW7YzxwIapOE+z71moux+W2XJsse8LX6jDJm3D
yrpSgupgL8NklyqoEM6pnUJit3ItIYzgECqUrv6hL1i1CjMlojpl7FMoELtKV28dFy1/0c9YthMg
6BQ+3ynRa/m7/2D4bHLga69UAUC+q1Zdma050UVYJLppcZ3r8hSlEeNnOqXhERLjmqlf0ev4EKHO
XmmTrNMkSEC1Nz4EgOMtQt6AM9fhihxpNQ7t6YMFybVc4BnUfzQ01ykpnCVKem6l2n9McGnUXaL+
6MuG63kYRDR/WDUC5k0EBbXFIPUSUL4tnHFIY/dAl2KtGpgTTZhBKnEDXU8YnRhgHkfHw4ZtFKGi
YuhmFwBUs8A6k79NZao8z5+GB09deUsvLXNEMvFnlh3o4yBd/oljhDm/p7admIlbmoflO4B51QEj
HfmRySBv8xld5HVJV/2KmI96yvzn28TAVgPnEmGGv/YCRe+sVormv1fEap+abEKggSX3L2p1sZpd
T3Wm2hf/Cj2yKke7rbXyVRp5Qkekq2FEZGEAOr8HRTQLMeJQZQCbP2OEBuIQAj2WSewzMDrSK6ks
27csbCP5E7V3G4k06To2HZfLIufMcADVie9VLThsMLZNe6saHkeWSNvtj0HnJaQk++U8navR0H0K
o8Bu1zmU+EkszUnpd70wqVIZL50St3uOAW4FQYveHqFsTDn3v5Vdp2IZ5IF4CzPPa4nhXYsDpS0Y
Ed64h+aEtp5encb+q2nqiCYplEkXyMlmqABfNsg0nTGQZXP7/TdNKb6tMYgUdy9crDSPzCR6R9LB
X0bSqd092KRVohFROtCpJBZOcfUIBCLtyDUqFMfKjKz60m3Ei/oF46nizpOseo6ah1/JB/KulR9j
xucdNI2qn7aK3oogEiy7UtzHOlUIoqQ6fzlOiDCvAQbsjP/peerSfaQWT03+6NKTQpeBOW+sLllB
NIHj9FOi+gGMdmH58IsUDqTQHRmip5+5Dkh3Uf7Qy2kGwbf2n9jEVJbptwXr0goyHLPdSML3xLY5
KUSCrXj5yPRB98qsBS7Y87dVkJ6+GeuTIcysx4Oo1ZnrB/La2TPzqunD4GU5oPGxepDfjzL1kg7Z
QjxT86H1ndvxryHTztdXoLkm4+dEWtb8pRJa2CDRocgBIIm7KqnvvQecbWK77qTQ9gQ16uboAC0f
TmC1P74tnzWzFYcKD3XyBnqGh5KOMGzOTOD286DekeE2lX+QuoX31N3BZAefjx2io7+DvH5ntlXj
zX8q59qUuf1g6bDZn955wI1yN6fQVCeRLWnnYVT6ufHN+J1UvzjQlTCmnBcpserfA3XCeE/nZn4W
et4BwlG9RNBxcal+c1cJkvOVxj3bJpU6t5ZHcN+KfAr+ewPCS/hC0q90OmTQ/GaIhCqQlGAwW/82
m4FvJRnomNULuVeYST1afgXbsmXo7gojwQ39ha2KuSURD7lyhSzkh/tGx/LYR8Lf0pAuMkDCNGzO
dNkuoFu5UfHt3o7n8XOsBRBZ6kYS/XhwFP5+pH1x+3Wnv8b633aHIn2nftf3XQFuCR4X/JklXq84
Sc7BNMwGaZyJqLr/48Xbpxg8TACj1Jbxgoo73f3XvWaPmTYD/Lb/JSzWQqA3scoAXxdpNlt8d40s
JfaJZ/xOpGydFk59gGRup/cuxH6OV6+ywp7E0l5HH+wkKu1nFnYrObtyuc8qgC021xfIlxSA4e4K
lgrizKRTb5nCa65EcSktrEGvpncldKWUlq8craYQIBdgvr5X6II0QUbjA4Ac0baiedAkUL+Bxy6G
r+T8FRFeH35u0UCbZBDwMKTz+9cDU+jtvQ0wZowRoWymZVnCm5JST+gYSnTU8dOb79a+yaEkZ6SF
99DvwMkLDbmIrhIJWVLxyVwum8t1Ef/0srolpizgJqwob2OkgBz2IAQ83nqGYh3ATgYQrONivKNL
jFPXk1B+UixkeMP14y+VuzD5u32688Ijle9HJvJpClfMhEmBxcxYCMVrMDpwpvDR8KYJrGnhVPP/
Y+hJXziPDiC8nVTCUOyp6WWrMVsZy3CxavqA8Idf/IEnSLYI6N/KLJqWgtIf5AmlkON4ChWpgb48
4qrtalrUaRSXJy6TfSRxmcYcdLRgmInxeEPBPp3tQwfxC40W6Y/RA2yEVDaej2H9i+xKV9Fy/rZ1
zOd5hdMd+404HE25jxxGqrmBRfRDe/Ret05nVocvXdKNiGJzCTITzyMe0YHf8m/9t1vH4NIteRe0
2wNz0QiGjCSzQjG6kmzGf+2Vz0rzYwbkfZ1OvhXLL1AgK+C7BpRQ6w5eEyvqbZ/BjExK7QbWI+qr
g3+/5k8WJf3K/vvmKzRbNxAABhUsWo6l7kYfKs9fX65rPz2Alvi/Dqk1ffo5+IP00S2XbNuEsHBj
xgb1IEusebORdWJLbA9uUgE/zuq+Le6c+9zdFcWCH6/nZlNHocD8AyfFZHZiz9VYdUCdnHth+aEy
eyiaKQGpbVRFZsKIO/CMPXOVWzXq3jQI8ITjloQ890l/VwsiVO0T0X5FHChlD4NZIajEZmY7cBtK
7ZvZALjpKbrAD4kpmzCuSr3q0Dav0hMWLhVBBaYq358z8LG8jVBpJMH6iFNig5+Ld9n2FCMFqCfj
PsTbLotGgTC8ISDZZyUIcPLdej+cqaxb6kNhJBoIxKQSl8TCk52Q5c62ppPfkGDCbIOBIRMAagYs
cBrq1vtMQKM5qidmE+hX751ClNqnoxYsnddBU4XHIQ9xB8TCVCg33Oq+qM2Z5TixgCoSxg0D18B2
LxqByZ/EtmzbsQCdsGrN0ZLFJJqiC0w7Iypn79Vb0BqGdDgVlURM4Vqp5eC0WT9SUKy3+hhKtai6
2SOkm+5mRPLrii+mCYpcKx+WzbwDfEIRGWqh9eHigTKqRcqoUDOvOadaBolPZdpVp0lgVa5HUOnY
4yMtgN1pKjF9cVoGhlSuA3Kn9PrbMXeJZ7vkKJXWaVtdekDGHIh4Zy/XiSVKKYD1VlJni8hkd4QB
Sey3qkjf0cfb8jjpr/qcV4f0dr5RL5YMDPMsHkSHwicVwrmc78IzH35QQao6IWm/rgE+4wHaOykR
WrdxJUn0R4F45Ondp9vIjg/NSiqmM6KTqUwqvR53EryYs4V7rO5/ICzS4NjsyxSHrrikMLaupoYk
8t0lT+v7H3z4bnvyESApeilPWmYqIubtGiFbKO+C70uoflcFHJgAwCX96BBKMtHuIZliTSFEFWVE
/Q/QaZ8Olrizsxar8HXZTr0tCjAyWXfKQ5DFsi+0XREyFfCpqv1sjuj7aSp8MXJIFRTEEAQElIHO
vnOnnX7gXTTqjLK/m+0ZDBFJbEY/EnO5pyMjiXgLl0TN4TYACvnbttBigPyOfM8DxZu+uDeoaqem
qxBv08lrDmFcPmh7OcMRqkPReMCJ03om6i0xbeysAK9y5+D8kN3tA9nvApQ4KiERGc4V8vZYqgk3
13XIhIV2wePnO1hhKBDtVIUOf/HRxHKCIL/AjMOyVke0/936rLk//wcPnArCA2NV4TD2IRge8bLn
/wjdWCH50KrXciHubkVARCQqGj+bkKZyCu8iBhIFeeRdN4JlYqiB+gueZr1v5lage9aIUvobXO2s
Ji+QaXauzLwjeJQriIS0uieMVPpmMbjh6XRLSKmXZJcntxHGBiggYluAfuFYaekmIUi+2/35v8wb
1BbJK1F0JkIEIVveM8+GH39ujcRrLJqF171woi5hUXZvnuKLEnNV6zlhJFbLgQIy7IHd04T7g4FZ
SvXzvQqTPmGu07F67/+cLaCJGn11GN3AL6ac42+E4MqJIjPrOphlOd60jSfjfiMt/3nW9S0t/+RN
QThANyDLpOz5a+LVtfK6Mx1FmEKStpwYXeuoTNHwmtTXGom9g9O/VKp4awaprov2yYB5Px1D4dBf
2fgbu6bQLmZKj0iKU4+lflxLW3ZN3AjnrCUI83bsulKqPrl6NWq29mZSDG5c3iraEd+286RE5Rxa
wYpBV/+JFlXASU0oUxNtWgNqO9L9m1at0mK7Hvcc/1iwskyp4OzUJZ+Youz8JzyYEIHi04Px0zJm
jIxLfdaD9do41+cMYivmzmbbAJyorParL3nL6JTvfbZyk43l27Zy8Go/rT+uvO4tSEKE39xm6n5j
m5jkzEhr7ppn/BP++lcpmVL0pezPKA/EihTkvzk5BiTdrozSxd2uFwOrlHsKD+TcEoK4kKM+yKT1
hZ7mMXyLqPpPMAOczlXOWMj5DzNxEomUlq9dMRkaBVsT7qvdg+y2CwL4n5sHF7Qfp3BVjsxBaQYq
N5wSIEdPpbD1H4BMEFdLdNOPnwBghU16SkxMyPjkmdtifM9B1rCkbirC21XSadARKZGggDvKO2f5
05KLlgQyrLGQWWZ8KMJs+sZWDLUUYvpJlVfLolF/zdTsczZ0dIFmEEekUiaTCAMfzFNfZAgJB62w
wkYoQ2xLiV1ik57RhtaD3Aetel685eBYT8HLYc6fxphL0fDfwYTo3vZI9sdmZy1SxqdVNgwYXVLV
1lvF7nECdUiiW1MBiwJukeib9gMRt7aulPIUGpW8kuzM7P8xPgdIotWiDczSevJgaprGdFPlzw18
AtVq0Qy7v6E5nHjvPjQ5qFGyUH+HO9Xyt2gM1ElaMdMw7I1UqKoH2KTRjTtGeTosWUKrYHF74sV+
3ebVB92AFodziaazJLYv1A+gTxv8mjISPfi4tURVMODKKVIbrGk8lDhPtbymD7C/5WcPYVehwRbF
z0mZ/AyFDEjzZVfe1J3mxh7sZA0D3vhT8on+0zbLPn5xNa5I5CFi4jBhYB7haln0dIcqvd9fsGz8
RVdZI+c20NRlOlw13K/UKON2xJsUvdESB/pQh7cAU4T64rOS0ZQC9mVjtOLuRseS5zXyaoPh1TVN
57HqT3JAUPNp7HQAcAMhLpXpc23rcdCz3gYVaAEe50n0QCLHaLq1XObSzjatrsim5eKMpoVtLkdI
zEvGBFagX/+QML1OIBxaGN7U2bqFK6MGq0a2zqPamshUZcdWxr0ldoCTZMWbaUHQIAOpAa3hqjSW
C/oZJUzN34pcNa673a9pmJJjE+lkpXUVnntuQnikwP2XXg6UB2C5NJ5EMq0Wg330p8NgWgB9uaoB
qcR+4QxLNh9OiYfgPB/HO783QH/y/fh7KlVvI5OHPIP6wt80ZjL4rnI+FXjmPA4waXoGYRvgbzaJ
HxC5TnBibR24+1vjYP+PminilU8YElLS3kZn+ZO76t13FEFsu7qpJ1oTxAU54hYvVUp8j6qtZm8g
Gcg6tR51VgVc0Bn0dw9zisgpbtLPutfkJIgMScOrpZBAFAUS8A7XKOoMyCDd1GTk+BtqxbeaRqbp
4KI8iHnKi/is6KziyJFJxMexrmcDeA0I04D/uDIqGEvQGZtVeV1+N5pe1BsRGgi0fDhXvk5Wc+4u
I/wGqXmHWQDDPRNFnIVXPPmRcgauUrw9gAuFYpWILVDc+6e0xL9D3ZKBo/aQj5kxmZmWKWqbg4+O
WnWo8HWgTzigKhrCi/frAcXgx51WBKplBWNq/A2fpHkGb0dzSvNd6R0+zozhVtUy7rYSUf6yIIsm
QdKDx3qg3fvB439B+5JLLCLcUo9orneQ5U24fPH67Tn+ORWMl0U7I1LAD8S4oG0+uSRVlTsm0Fsg
1vnETmak6fKqtksKeTDriYvIWwFeQVW0JC8anzw6GKHaMZClHL4jMYmm+p3zRsFnJHr8Mt+PnBoh
7sFW8nUggfpDN+KC2xOYwspQFE4hOU3795rhj+n/rp6TrC1qgC3sJv7VP72Z+JN9V/yCZ3u7Q8cL
PzW94PIQLfKr7MxgOQew6XwWe3Kaz/aZFjOyto0w+PNLEPdgLdSAStIG9BhgeAe0PVCrwEJWyiaZ
rMjvM+jGnTWG0ETkDDHF+inGQEoLe8bDMbUouUqHEo7Ulr2L9qgTlGrgTKY8koEeVI+hXqDT0noe
8+Tfs3JitXwm3lmpyjR1RFledQQicbtwnz1e6y0xBGxs5VKcVK9KVd68p1scRTuA394uUzAytkEq
f7SGVcEpICXXCBxjGkrfjE2dOibUO2IvBkL/jIRDS9rPVw58uuCM6Okpio8o7fSdxSet0osFXeNJ
3eKJ4TUmTA6d7fh9UXS8R+Cvpj7bJlxfEN2PIxtdqLqFOtrqZK1Pp2GfPPgc57KvwAtj1tNZ1yjv
eixAsHtYiW/TFJU/ABXZEFVgOAKLZRdM1ix2dsPqILQdMpaszYd86PzesTqSFiG9L6zIIEqAPeX6
tk3vxBj0bafl/7rElMNNn3MoGOCoRYJsmocSagb+DAiOHqSV57D9OrpSLaoHf/VR23P9rgBod46X
6aYgU4TL4AFN6UEXUCriI26cA6pVQJXU+Z/19Bc9EX1HTkBgEZ/3612nB7Mwt2qr/HKdpmbvj3/R
9gyiamzyC3nEj4nvZ9JR2te+AS0o9oA2znyFoOYa25EDNB5UuPmzHlExJ7rqpO4jKoedkSXTrW0e
6shulsvT2t7jC5sSAkT4hAKzIWH77GlpyUDAEIAJWbxjJtlU3E240DCu9KSGxFPYl4sX6+17+0Fo
Z8bq2mycgkGYUbCIewB/K+L9xF2goIGtJaFBQV06Weadn2Ft1SiO9kHkcwyBEsdfE/gn9FVGZROe
N02/IE2IeaAswl3zB09xheg14x5ZYCeWsXUrtIl3cX7AzYsJcM6ewezkiWgZjxHKrOFZuwlClnRM
8kYPoKDqZS9og/WMSyEPapdzcHUFnfZW+5dhzmnF4vvjQuGeqqbXHP4vyA8asqaxL+QBu0+1VBmW
/mAIxXq+SXOeCOcu2gtG8AldTHJcZumUKu5vqyzrLvxjtjdDkM+HjvUhdLMzcd9STSr1S+cu5EWg
SgpM7ljI1pwG2VIwSfF6G1AbE5x26y0UffCanMrfFSlDxCT3nn8ECV6WtUPHWXqVqVptP2wzxCzn
yK7/JwtdpdFrsseEZHnDTnQxoXnxkxvbgvMHWXW3DSYfbFIcEE6iZW9yERgc01SfaoPdvw9aIPJk
dvFGwVz8QHEjlWpT9sPEE9b+vyVn4FQvkTSHFTTeOXPXTujFWoGiQVUe904/iSqUhiHqRUHK5v2+
eXwAoRhBPCvHPdwAwX8NAMRfrakSZaNwuiR3HMbi6QH9n5YHwI4kWwpzFYCTW5Flkezq5uZzMNU4
wvbnoyEYA9J6/WSNiKrlrIIawYMEQPDrtMa4pAjntX+DHVNBrUmcG9CwgPnn7Tb1LUVGMPxvBB1u
mXYaJdb9jpnDlIb5W2rUVytm3+XkptNlZLtcHNc1IiRimPozmn07e6+/SfeJhUThsrPeBd/wDyO6
cLrSy/P/AVpK9F29c/2c27YlUkFHFOYGAIai4bgcftKpR3xf+jnQQK+h1SlQtFMg5o/XumxTOLuk
3LwxQa5yhZ4eJIfyB1sbWSYL4XaNTZDInsVBf1bWpMJMTMYV3GSB63krhyXoMjT0OzyRMd9DL8xm
px3NdnAEEIP3HaRpHlr1xVFyraZ+apSAVqUG1tWc88586AfI9tpQfYkrSFFQtp/0cgwIbONXzxUX
UbH6rY8v7XAPpwd/yBmMVkflMYzKpvhTrQSJWHy4vQNwtGECim499qz8uA5dApn12P/QKpM/p5Ly
hvrwzsrYTu5K906YxfNMz29TJgVV8iCEa1oBeWvwvBZE9oxyqXqD+HfSBKeztVT+d5Feam4fb4Og
JNEiB/bpEwOmBrug65OXcnyNFtJZdiJHxF9bURhzta84EhIcX+8lC4bRg1iglEcb+YgOz7ZvmuJL
CbLR5oYRLlAlwBTYAS002j2JvXFHBbzsMTRnMqDTX8t45TLzAyFlNnZATzBUAsL0JxygkdnzLAQ9
Gph2JSnfGM6b3N1T5rAG9Pij0XepCaPKpepbpPFg7LneKhEAOfE/uX3YQdA7Sci5nNRD9oH8vW/X
EM0vapO/8cYNhE5H4LbrpXiejfLcVLTw54X1G8c5iKIghRECvuTuR+lB7fMcsjIfR2d19uhhPK9a
uT/eYrdtV4twcL5ghNVtWk1MPPIql2QA+F0sLO2vKyLG/Alsf9wumigBBBeHZacXeddrOIaebHrK
xvg43eR87LV9VvF7c73VnxrQ/BlmsGDooosOkkShQG1tnua8aohEST8VVB/olo5QJl+EGLp3qtm7
FXAWn4W2oTLYw6kH8BV5kyDAxCPb1vuDotSv+rvahbbPWNdz7rxPqTqduUw2s8fhiB4b55Y0Y/Hc
zaDdGoZlfqYAw1gPZ/SyQFJfCeOSRq/6ET6EkL3EHj7CM9HS1y6T1NDrc+5TeCGLqYmtGERjPk2c
P+MeABI7eK8T0MwYkbB3CHWd/ha4YFOp9lbm0QX2M1NctBrWtqM/VbEXecpFcQ11EhTeAR9bcMvu
6d7k0qxYYJ602egZyJWgrgBGAs7siGQFtEVOrh+GLjnYUJ/KHRNi6YY3jBeR8dQ9r56i2d/JqAYd
MnD6WU0dEPKfbvZ3nfWG6WkI463Xk0PYIWvzKqFAzOGoHU0B395cVcmdkfbMrfeGJ3kN/1tmpb45
OewA5AmqDQPs7iBpAASME1xe/DX6hf0+M2TSa2eG/xwEpIy18xvCyY+BWXEhSJwbgxHyN49bnotE
OKu4Xhm2Fk4GJC+nR0O/JBG5JtQ8wM/qiEE2cGk6mvoZRRXmOEAxRMNBt+gyKqZJulupYSaWY0Wp
dY1oHPT46kXQiILdD/eaMw2fazUZPr569Wo2EfdYLSk/Fc5gUn78SuwhIixMCmCmgkHVwNDLfxAu
dbt51dDwQHHyi5Bgbs8OVW9ks8JPTpnit/kbF5JmUwRRMLRCw2kLQ6KJaW9eiLnbEpShZQFYe1ew
A9KEX/D7F8VqTZYGonKk99PEulbB4f44cZ8VsBVSeTteYdg7I+b92WHCdPeFEXZY7bncXLB7veOZ
asOfng1i4BSJ0qLAA9ynJ51AtiKxqN+T1JROU4yRzTLgAUYAEWqR3RsgNH4XKGVd8aGM823aD6LQ
pwXmV7wkViUDF/o74dfbzsuklcONOyXTo7VE9bldLsxLeGDRejmxZ04LIlmhk/Igf0aGSLK1sk8j
uZryCArTp9JfmL5MEmlPKCm4wvvwIT9vVPhmQSwIIcMSCfKnR3WDVMHWZ70RZC7EQA456fFQf8Df
UKgw/2oqyzZbl/Shfutkqy3N2AvYPWnbmBpXunm+33xbm3oJ/bhrct8jxqj2N7qCVcpqtkbv8LL0
fRq93cO8R+eYcGgX5av/j8aIMnOsbwjUoQOxjqoPaMyDtbCnP4FNy/Hi6Srg/rW4JsmUV9hpgtY/
+Yb0b6dq11W815y+ZERQr66E1+pCg3RHs61YU6VOZLz6cN76pX/4dCj/AYf6Z1PpezHKsQ07lrQR
SxzDwZeaU6TsoTvsTTYuP9KPCXcIersuHiC6YQ4dx52DddTTV12BmorTigpVwFEzJxtxjii69jFD
VB/XwGBnONuDAjhy09o079EGj/UoELoULTNnjEkvdXCCzAcLq6HjqThMFqN3YqfPsHGL21kzFM0w
6C+587jdP5Z2ThsPCo37doK9U9JnwbNFdVMVQGEJ0jg6bNEl2jPCe7Q9MMcAXT8+4x2WQZOtwAG7
nf0x41Vd+6H/KX+R7154QpH/7X5cZAUMbn51gRIBOy7H+qrqJCGefjBcmqRKjjMcB6Rp7Ni48sI5
siV+AMAEORYShH/niwhoXhlekL+8A15nVUBxyj1H21HXXZf4iTtlayyZrBoZRmwPc0xE6lFaRklF
s2YUgK3+bxQtT0Dn4olwT7kkQyr6HSwA2Gl+kvFlvaChfBq+TiJXU6uEbdo98sb3F92NBY2zc3pS
HKEMxPivxgSLME/0KZapoUX6Oi9xbx36WWFA/gMHYr6fW/G+oFdoMtwVkicrT1ckB6Ac5TrvBUHx
zY/g88ExEGrIg6F/DUpkTXDCQiDAU234aiwcDNlifi2NCWEZE9jmAoMtOJNbXTaAK8djAO+jr1E5
3AvAcEun6zBUAZwYHxOPyxCiW3jv2Qtqrc/j4Nc1VhmyHhkBmsEVh4zn3cXSF98lSQQuJL9uaIaX
3zJrt9PhdDnOxZEhAYL77ajFoPt3ZhWnoq0uXTwjurgRlbVcEJB4eEGGCBUQJrF+va83if136FVc
sKXUPPTdZ2kla7gyFjfv0GHOZXN/cEOJf5cJLPrtC+vnlscdSYSRzVmYKXNDxQefW4cn3RHF5Yda
Ec5jGgxdmhrNQZWBZq/Ofw0UPAqugXI27zw98/Ti+bGx+6xVei7U9+a0RYl6G+7TFhG8dwO/eriQ
cdKJVC/uTeBFpx6qCWnRpl4mdM52BEtvwC/ggk71yluvBtuyx8zObg5LKqLihBSmFK8kIAfob/Im
4QO6FSc0Mp9s0U0rp5LOe1uYYc76t/IlwqL8vfmMNvrr2Lu5fxYF6fW+5NE6hNykMJv0EL47p4SC
j7OlCDulc7EAfBTZ130dE2YW4mod8zcUUtB2pfptG5SDvfpuRvl7EMcQpAyD2BpZ0bUflqJCBhiQ
SMxCGo0CKM/Th0EJUTJ3rndRjWNAEFJaUPnGwcf+pIVTotXhEnTY5XYyMx4bDNXZL0bQTQqhcNtF
WakGWstK4ibkRVZm4nEGHMXmmnvM8GKpBNz6QjjWi3fWhOQmiFjESgPE2AZUvnic7MzskbarSSg+
vXyi6kVgIw+Ii7m5H6uNXpbOnuazUMm1A2LEX4kzWvKBAESK3XL6goRODKwOrA+TIh+vJS3TB+4x
rNi7D+u+mw9bPvQONWVxs/lozRbS0Mbg3scC9Q2yshB1GAX8KFBsWMVCliqKgzSIGBkTLZmNx0cz
GOMZfg1U1n4LJcFbQOKxRXJFeVcTmlXn6ZrSS6OUN3yL/ObI9RtEkUS+0NU6NJsP54QAVHS7ywLf
e4E/0ZVMQJyN61Rwt4olAstEB5XG0chEdO245pBkxigeE0xlt5ia92gdoGIHejQyY2MYDg4fIyyH
4d1tJ8BocPstnP16AfFMGWMKJ5hvZd2nRkxv89Othn8ledMg2Ev2dYT/9f516Zwh2OYAcJC5rUHp
b7SZLB3B4hlUs8vrj3ZafXx/hh9HdqFgJigF7Ylpa0VS4o2PWTSyVaLPQOtorooTgcFdfbNkkHja
7KJ4CVHeczxLlS1jxh3+wZ3Hl4iK5ci2JTZMuPmtQOJfIDLH0O8pKxEBgbLqHVZLl7VgljyzKV7F
muA2brWCaG+me5zzdS63qAB3oBW1eGOmyyh6x0wAJxHCc7X8O0H38rt5A/8a4qdHdIdkfwyXlMsG
d60Alk9d9cAViV+f0EuDlUXWXgas/KtXeStwGRIFwwvAQ0gs/H/EIVSerFgmKl+qR8WwcNqrCiVe
1J6ZTKxV/PkEYbuL/Lj5t7uJdjfyQwPut+GkX80ejg5CkE7NHqvZU1cOSw7pztEtyTGClrOqSBmg
yW1faY5xNbVaRhd8U8JN5ezCviN/KveC5sjuny5fs+stXsRkfdmHh6dkskdEKr/cSPa47bxG35Fr
WrjwsklWQRf/MzORAu/Wyd6zROak1mP0MohoO6fHnszGXlagsWKRw6/MBwUAf9DuYMQctakOTokk
azP3f1s57FmQQO++PqtEroY92feCn6nRnGcxoyrgyD1YYDo/WQdTxUSl/rJ0jCH/ubv3SKR+4toU
xjXQzkegb4JvoWG0mtgvjeKUfi0ATyZf+f01S5kQs9gPKSs+qqqrVSLPjAxQC19VY0haRtOlZvkB
xk8vhOPTiZA78jZnKv5CWN2+fMaM/yAF8ufErojTCiUba/zk7T4sv4fqzBYOgpNV8HcdqzI3ruJi
8iZkVlkJ+Qo4uDryj9OuSRAmMaj9xW9usMafMgBlEn+C5llo+yJ/79eOXEJSOfoE7TOjPMz+BHCF
ynKierP7cp1An4cgG6epseuXx80aXtQazgnaaVohtw80IIMYZ1U2UHVN9QuGc+jS4i2AOBvDMOqE
mOVaWqaujZbMJxyGEw4upML9658z62qg4PCgwFkIvj3g4L6CG3rJiBjBCUnAJpvyMHxL/zMh8I+W
a2MZ0/kiLlRvYtaal30VgXoCWWfUtpt/znFSFFz6JMAwb+wo41xf9nhH+T82B5NDKqVJbi6l7tbN
kwIQsMFkeHtyiojG1AF52cLpAMnSxdHtYej4l5eZrW1KtJPJ+ULgQy/PAvtzxkLJFUUxWTuucELl
fbcMz0867b90i0QiTIzhIDK/72Cp9ecGqWqgNkZp2g3pNf08wpLCIEa+q828QCKvmra0B4LNKwwc
JNpkjIQHMQC9yLCFVtE/NYVcmdnkd+lrAfZuC5MDx6UKIJXJ7sPsfk+J4uG2bSnuqDiHWKsPaYzR
W3dntPm3F6LKqRMpzOym/5nxXshA6tVmcW6A5SXc8nJznRMKfAdWG/I7rVfLj7S+BNJuUbQnIEgK
yRrimI8AHdqmSYMAmyzeX5MDmD6clzQsaQXRAmjJGjax1fKQAzUiC8XM6fUpdHTgldMnmvFzF/0Z
Aj24KKJ8xtfo4yac7al3xumd5ehCWak2XiuZREyASIiobLSpY5zpmFGPGzUfpKALQayZDLgOmZIL
vmrxcIcLl2n4CFf5DShzmh2FQqmsbv3NnCWrM3I0PV0XgO7DERPT/IMbotmyrosIROlpI+1LOSyx
ofGMCY3krH/0D35cD5nI0KHIZo2klPoLSSf5cQSfarnZJ618gFWxcF2W9lQIPAtUxjvFwil7QwGo
CbKbuLad5zGPG/68WLYglJfrz61jdP7i7iyQOvQ55r55PotJ/xxEzGpBMIPIYX6DlBfFO0BeuFBz
vl6o2ybgEuMQyFuxEoHFth1bYB6dls0yzDvR1hO3ODkt4Nq4RtoEtnvKC+vXlhZYWx+S5ksBNo48
VaXIXuWWYAIpx07m6wjcotZ0Ln6oF+db+BEqgHi/BI9ZxKEEATwyf7twREtOyS+KsPLKkWDscjxO
UXZ0z8wD0X8YtGNSgEX1lCwOYLLfo3V+JYf7ZjJckK3JWesenPM6tK+bPcX6miptYKoM2mhbQf70
Dvg7heFIWUdCOykwLkadLQ7K858LR+DDeC3HXjIAGveBQciRX6x5Z4TWjRvk6vzDF72Na5jGJuIS
2VY4xMAdjeHH7eFAbPHFb7A57z5YnG5kYDaqWx3KAk90frhVr5LV8QhdOWrA1GG45X0hXczvEsvX
8pfQWhZCs8p6ZXkFD0wOUTj/cls3d0qV3/FaQgwSwUMeUo4XqyA8uITeFmWO/eCbdZH7c8XsJEQJ
2VUAMrzZL+0ABg9NLrr0XSmukNnMM5rZQgF+JKZVPRP2PjnO3h3I1GdkDGxDK+7wiKVsfSxzkRp4
VWtrv7qLipvlVhaWyPjZY9RN2YEBfWtyMhn0AM51GI+wRQSVYgx/8eXkJzhPCEOk/tJm3ti+cZEI
ItIhOv+HayI+lDyztuWK0GMxFfVoHA06r7OHJpFpGn6mDqvLDx4xmR2EtUdPXDCoTmPmEOkaUAml
8H9R7ShXJju0Z3Gp1OjTNrf2keLDUQTxXVVFJ+89RRbyp06l7vfTxY3rFu9tU6HHZHGoY/IfqDcH
KIPiwG1dbsspyVb2InU1TRhp17En3LaXwqr+b6IiPW1dlKvEzszYfM7kfS6Z6VMQONd1JCTRK71v
J3a6+Nr0UNyA51PAQ7nHD+fcUONTon6/pOytz+6xVdvKXsLDV8XG+eMde0ElqXA1sbDwzMF5U/jx
wowO5ZvRGrEpvkKOvp84BoZihyxfR3ExoNb7Fuel8O7xLdgyq2vqXBZREell6YCgbZXO/yMk4ZJZ
ltQEOR9jbvgRbwbrY+iPWdS2g50RYnT3yMG6VQJDCJfyldW1vhY4Fr+Tm6jyFrPBD6nl6JSq2o4T
qihxIqcwBVXqEQYuHev15utjlGiQKaiXKgkTG/612f7dq1emtDYmzxz/SkWYa2Hb3YFA1vnKfheJ
rTbTO7Boi4/BXt/w0wXcmcQENb6c/jZiTB6mIZp/EAmR4GO24Xc1BXYEIAZPFm4XX7kUEeVkEj95
1/f4NrVs0Rv3+FLGrqa+g3bk0ylnyA1RvvfkGeFvgMg9qdsWm2AG0u+j2XouwTI925/T5/M/vwiS
qEtCgsG4XV+5zbcR1GyX7Gk/c1Mp06fiP41bR7fPLnxLbHFkqw94Tn48ZC5iTUwgwlR+GP0QC4NZ
Xti4LS5Azx52Q/FegFSWw5p4bMTCJ4FtsVCEgob4vDQT7zSqO3v88Ih7d6zn7wlujNqCl9v84TvO
Ak8bLmroguprsZebkqgykWdoy7pxDI9Ulvf0A8LLRAaJd9+f0j6ZF+Dxq50n73CMMnkrPPG+or2x
RzVhNTdJDmxWBoOfOYs6uadBzvS120z3Pw8ixOzndRh4JCKS9XN/pD4mDcFi9y78k1amkx6f/yCr
ANOY7Tv+LuIrVo9hYxsDZouf2kPBFJ30YNf6DORTslhUfnEIJoIqVCaBveWcfz3bWjUxcl7130uf
8V75Q8OOkCzgYZszrVq9VytWvndv2TFLDX3p0dnu/3gQ27yDvQkTc3IrWJaQbH4OHg22mOps40rU
qf8Q3IJf4yQw9aNm01sitHJNaXHNPglx7CGYVbo2azsp991yZCeecFnkc8PfGYjYv7jcXSUaS7b1
PolslrEnHsmPi4nV1KHGKztQFWRmFzshAkbQMJ7foUxQr5YWEkubT1EhP6XIUhZ0sxNS4J04SXfi
YRE4qa+3wX0cthc+xys+k2PONOUL3AQoEZ665T5So6CE51k1+uvHggIt0G8Z7C5IFdoyt42QoT4B
2vaLjcXIEriN8TkrZqS0eZRyFIw0cZOdV70obnjInxCeUmIfBH9GmE7Sfx1K7Moza2VvHwQx2JpB
IBwL+7iB+YgxYO2zvQ5Igalez/kpgPHEcjlwlNyTqR9s8/bZzHDJANfwFqyYRDf31+OGmiZUvBYl
i8Ef69SRLbf5Zw4uCxVj1TdRCfmkugspyXD9NXp1DqGbneDfkWdb6Ksg1RRMCjZGE+713x8Dr5Hf
Gd6ZYyJyzVw3w7IkRxfnIOTrcSuF5t0wrCtK+knlccsBbDZN1/KTtidvuwpQtHgvLfjCExi1nqU+
7xDEzJrpmJOwc+KrlDi5uFGxbhBG4aHCdDf3QW94If7w5hMONDrZbWQ4yZLy6DHTDG8OaYCMmk+j
xhpEkDEaNU5opi+vpSBYL8gYnnZOOtgeVBpfHFRLQRBwhtK5SDn+7Y3rFGzotAOHvn6qdci8t5KG
tJe2IKiOLfAo7jZYZJXc4G6PXlxy8S/acEQ9/1x9fAF6XYNEZb3gQIwvlz3aRAvvF+E7oMx/xZMb
Fx+VUj49XzpOb9bigue5LHBC7TiBd+d5ZXbjWOH/hmQ1zXYcDCRdgMWPfuVxS6JLZnItCBcGAdqQ
1TUQ+D2xy1lYwHQ6w/ojMY/8CIHug6AIGh6nFtrDdBgihXcv10RKUE2e6kbWjwhUE7aNh9mmtI+l
DZdcx6FM17IOglvtk5YFr+ZRMGxOKHNKY10iEmzerxhl8FHzyif2O57pPsffxM7wAdeNo31eVyU/
IVQcvq9Od8j+nayUuRIlm/h+g8wGkjl7R+avDzXYqRyP+NQfTTSrnvaNweie+ajDHgZ7TJ6LkwNB
TLmzTEOZ+Bl1PQJSLSEgG/pBXxs5Us0ibgJway3ag7+ehqZwgSD9YDse6cGxnNK6VZYtwIHqN+wV
lmL03vYcK9plPMh31lxqScVxYlAJtjowbs52LfZ+RMWaF9duzohw+UeIc5/A6dqUqWsAmGp84X35
87byTdRqnL4BkTVhwJTYuPnz40WBJQsrvriS9xK1a0gZejTGor/5U5TwQfV3OMoprGjmo3l8y7Ik
+35jn3oy2j+laz3UEVlXKdrLRMBwZkV9JZGaold980SimL1LxTcaJnMnBXwj95K3XKZv2ndirTG3
DRNMKRFZ3/5prZn60whiIDJ0jQCRnbFyxMQuigKKxm4uVuOv08nghs1PiwxDL3sDUhlSgPBCWKH9
sjDJeSxiycqvcBHYe0vsRVd+OZ8FDUI02vu8M+BrjWidiEdv9iNEasJGRhVLBcnYxgmylrRjQM3d
XobjwYdvkxon9f6zJ/UlTmouVA2L6NuP+fYJFOviyhZ0lcp8FqKnHVge6ENnQekxH6zYXrNs/mpm
ciTLKiisPYStCnrNhYsy/Lx3zG2QVrDHYj/CQ8wwFrkep63c9ha1i90reEhPjV8qmOiN0Fr6PmuJ
QtgoUeUmgd5ZNi3/kFhTsLSXJa0KZMtk75SMwhPYtaBzCVOymWT0pILAa5s3hQRVzwXBuUL/hc7l
eR2HuHIAxXS6yGUM9kA1p76dr//mlpfTvnIXWpgGJWnrJXmUIDqO/U8m9TeOhqwmJLp1uDamPI40
Xry2+qAo7Ok/yhepfnLfkSy5138tlyoLDpRsp7lQLyaGDKP5JaSf8TZg/Cf7d/5B4U2Qj+DmZXfX
ikZ/m9ZCP9rtjLSgrn/mXiP09JyqIkJN8nmNHs9IWNvq8IdCY3wSys2+GHH02e3XKOuJjtzuAHnp
RePnJsqAWCLZD6x4bQPGl8btGnMPcoVogimi3Pgel4vEPY2iKIBaHrkhVMVZ1TAM3SqftsXJmWr0
WNOyeMqUrOsUyyFeIuPfB5Xt1Jba/wU4bTTYcqZ2f6f3a9/Vb6i4lNCfiuRVjN8/a3gSRvdFMaxG
K+cj++jpkuxAk5gjl+5Vmkiq14wcMiJozMSgZ3yZHQNpU/dT5JMjbwh4cFhiQ8U+2231HzuHtoyD
2yVVB/xRkFURQWOuhDkwW1fTb4Xcsmsz6QAKYAzUezSfyw4rumxWud637M9IQ9ozn0tC6I8XZPpc
3mR/5W5hRvTRpUJsceT4M8F7D/Q+FvdOWvHSxY53LddhUg6fODdhaUSEDSApO/QUHII+RSR2+CNT
RUY6RXP7aMFa6Ndl5u5H7B9No4IpbxVIQ+Evv5lqnWsIH1pu0kmxW/X/tiAp3LSKRTPp1UlALt+w
p6nQqRXvEpACZYzvjlN8YYLGUfHEcnOPlCNdCIgv9/1xsOVKwbvpWb9rlSIEtY81eThtQtQ5ffa6
zJjsN6yr62xhy/gc61y7DSu3wt4kr8Rx/BCxc181QAuhayF/yVPo1+YiG2mwR5cpyHOIYI/zFxF9
JZIz0lWxqA/ES7XCyJyqsOfKoyQiv9ZrL13+ojFkGAhXi751IGu09guwmf1+hBlMaH4vCCUW8Cho
VV969ekCrw9K79MBKg5R4+7GzXQM2zAvy0TaRMueM5pOUgygZrYluImGIRibQ3qDJNqHE/skjxVy
otb1Lb4x5laGp56SLBSdNzeB4c95soi7mgVEOkVky+x061QfT4LYCJpDnAvIG8+ujNtuTavfEFhT
Arfxg2KYjkaNOHA92UBPJMLiy5UM4KGBreWMwFOD/HMqHayqeSBZUZYzryk/4RYr94HU3nVh/w9X
gPJ2al0DEaJFZj69/ZjgVPiKTV/9wuhJLxsMb+fPGSyMttc++FbVh9vTJRHQJ0fBusTcNMg5Xeor
ocoH63Zbmf1C/UgUbMF0A630WxUpUXmFi/IFKyo4rRzrelnLqL8A5cUflCiWDM4pQ0KOijdtlV93
ruezcl9H8QnYzAPBfSDvVgSLsvJ3jiRILa4X4F31e01qjHbnR3cZgUYY35UcD1vkVDrnCA/CHM3A
UN8LtIJGGNX8J4wYvx+Kt5/HJLKrM2tNOJH76pMtgSlnsvSa2PrTdOt8CU3KxnrcwKTUADbsS0Bc
RC/elNy3d9qaqRo0lR90uGwLLuJiUECVXEqqIfyegDdto8b81l00mZj1QRCfolqCD3nJuLpUlewj
nBE+CJjzHWer5oqo33TigKMdwRnt2VuH7LjCSQB91nXCNYeKkwNWheGUOAhmqkHE1obrT5sO5ubj
LSBOtomuxJUKssl2Q4DuCaYRKdBrWMPLtHKA8+hYR2fs2WRoC7N5R2ri9fLVYbdn5HeGfh66Wncc
Z02LP0VL1jExVyxyjruuZNTPBUXW6p2W4txNJ0uflgiI2qhnjtjZ++6fnyeXtiYx/RtzJZbR+JrC
HE3+21EBdM//SCSeHUI3TYMe/fYFOR7rzhEK++EfAEeMvyJfccEEbEj8fQL/BAe7qEHMY/1ueEFz
gqMkRoCHXL8XDooPa0uOKmQgeO60XVGHPOEONkvXKA7xQyjtsHXIWBk81ZaogIHaXGe/7r1LP60L
b7LvYd+6CmWxMi1yW9kYuNSmxrHiVA6Fx7oW95Y+jZIAtWX8kcfGKWCa8Nu8W5aDMt+RZqaAxSvH
cmJKnVSi8EgzoSwuZ8Cw1QmH59RiEBh2u1oz8pWNEPnX9uZ/Y6eiJI+ah0uYmtDETgT9EhvoaUqq
XPpDnocRZy/3kJ5MnvsCAkc8xyKlggQSxnAS2UpTcfMMsCeSIYyzYp7bccYz8IkwjHGKpDWvH7aH
kfqWiqZzb3ctvgPaWGa9zmA6/O9YZIe1IfMf6YuFr6ObAfDOF+c0YUTjL311e/4VYm/ZZzf5jyk8
y/+zvi8FqeSZis/qAiik3Rhp4r/s470BJwhqqfIYBPczJ4EcCKutUfr4XXrNnBoUVSYLRHAdPxq4
5MGjGbpnL/kiUzJysKqihgIxsVz1t6H/wjZaPlR49U0odDSNjJLceFoRzFZtVzTtjgW3JfGCSsW6
2CDZfHl5BbSWYm8QllAbSXs+3arzMluO1/uAX43n4oOb7le6csamUbf3u5esOauPoYOwYyDFNfgM
b4rnvH+2J0/atgfxsu55A32AlxQbnXLEXM6dQH1W2ne9lh8E5P6udZ3xuT+i9pakKuMC8yticxVQ
tzljUSyrQwG+XWpQUY9xJ6jjX6emng2eVVnwmnJdW/01lyl/s2fkCdZi+MlGAB7e2ZcDlf5GCzeX
UtCeZHOghVKzdqtJdikeCZe3etvqYq5vt4AwUZIuX81/Z6A0d2/5DThe5ynfabjJ/75KYnCEg4oJ
fVx/ofisnFPZ12vRJYR8h5SFvRuCm70BT0CMDQjGwB51oW7v8vx+pnU/qeiZ/ZDED1Yo7U0scK+9
IH0MlZOph5l74qErs+k2AVFa+Pp37wtjdCFOvxAfS8QE88+P/rMkUuvtNm3VH0kqtPGqFQ5AZIdB
4jP1gQiFXAnqfT4de4QxU4D/kDlqPcwb10zsh3w7z/0ZqLDL+AHFdsX6djFcZfMxugIv2c1TIC1p
7wUc6TJqmCd9ShM/vcDC9Ntgyx7yuCHOQbN9fuwouNavCRcBN1cAmKSo0KBQqkxWrbCj0DOnExoP
9jCPcwxzXWXMsOab26v3zoqwzdSOkq8F3WgDmhhzzAF0He1MUUY/eLcckpSDcdp+g69YrP/C8lpc
dOjYKTy80Zp7g+nr9cmHQ7GAEOv2n/EKoIuSPsF2VvWoDAgOWU+wvSXWO5ebRc+FnWO4e37OMxW0
IDfta86efWGQfSe5dtHWipwPKx5KBNAHmK6Tju3zuOCxdp53Mgh6LGcoOMGMB8Jh65Tb3hKs1kxf
65C/2ktq+9siXzxr2EdtBHmsHNhe0HQzhJvl6HNbQZkb2TuQiM+UYvc2cN972tFxMq3Sqfkre2JV
fqC2lD2bD90fIBHoHG6SxXVcRvVsr/W0MiaEGUmA5THO2IvrIn1EyO+NlgpAEDujmQJMsmZN0lr2
KHh+IbAVqVZG5xl19dbJnAK2As47CMi85InNzR6EijkKuNXAHrcMpm/W/DJFRLEYaTIlWlsKLONK
0hHgcAsu7gs/AHTTY8XNYmqh73VfQ+6mK8qoc8wvOS61Y9cTslWHe5I3rMFcbp9RyGEXEK8p7M4U
aYybCZlGesmuwUSh3TEmHuyVd4AUScy2FHTCUssoOxpqWaOfik+Woh6snYkJGF8id/z8IjeK/P8U
qNI+O8Nm3kFmaovqs3OKfgFZ3zWYUMKBSPG8bCU2xBv9dprz55qg19TCnLtV812TkP1YiIvAlbZN
5pFhYrLORY2sLPZqwfpemvGo5r7+YbNqZqlsgMOc4TKIliUPxwuqxZdhzDmRGxQKk1PIDp4XLsZC
gAstg2eF+Za8FkZizoU+18BMDVWGV3jbUywfRt7daQJJm/l6wl/XJvy69CYM3e5hD/+aoZVadvQI
ndx3wvp/3drvR70+GbgHz6XtSitRqVKOxG9S+d2UStZhPpYKN/tUwFkGZ/Oe79IQFXByj7UfCU7K
zrhQ9tC2nEDEiEK/bjxrc0slfLFmP3sLv3Gq55uXL3u0iMBfhjPCK63K8WFX13Kitwf+IuIZohw3
m9gu8Pr3Gw3sM163uX9+p9VdjEWJMv2RDjBKWQORSb6YoQGbt7Yzn0wFPUUumkAvCgcU3unIm/Fq
gx3S/80r4MZgmpLihebShPoeP/WA13TIOaZK3+QgQhAw6DyFcORFgjwSniP6R43eOCFIxEIoUqOl
f8HL6flsUofBo59BAG34I+EPTtGCS9COvBT4aJbK1mmajTxw/foPgtFiGf158tRyS0h0BrgFYLoa
UpRWuFV7p0sGvN8UUdqM5Chj7dyCQru+EPaGppqTXWgWIqzPoqB3Dnb94Hl0eStCGvCscO1WCEwq
OklHe2n1Ln/mAfYUDVzuK/+QFyf6kFKtp42OANrpdrk1QNyw2gf38c2zoh9EO8pR2neoZ/4GPTGp
SPZKRPZg52TorQaXV8mW2H/suKVvBgo3AbVl+/LgWJtl+4rOUTzv2vpzxvllUcxPb8+ZLryMnJ6p
irBbfYsWsvwD0C0vJ+K9RLQGw+TPk5DKlH1bd6gSUHra11QjngmqhyIFZxMFSLjz8NZD3cvi43Tk
KlRBPFgUKwQoGvICGkx9x2QntBzQ3gFyrumpc9jDx2VCSRXw+qOrmbdQpTSydUR+ERcdRzuFVJoZ
DaFgx2zMzrk93GNwkUBvPNrmJvVvEpBi2LU5xrbiqwqvKhqvBewyozYdbspABNX9nOcIM8CdbQI7
3M8ZqJQSgC/lGlmjEQC5QSHK4+Be0O0ZPzepGTADF3+K1HSHXGIwdqmRrAfOiFp63fkO9Jrm0MVb
QQy56Byk04PVxNc+MMepyJWlRxO0WqS/UKK1xABNeMKjd1F94UzIl42JopfmLwlAAUEN1zae8+6I
1SZUWNbfsrHUF/uPz6QsZSBkgF0vfAt0rR/X/7X+2BFcY1hSfwAvfkOUc1UYgM3ESH9S/ujOpOjd
MPDiW45BSALrNuCSmtQCxEI5sw0noMXO0QUAvM30ytOS+T1vPW7/U4VKFDDFWs7nU+bnunwz1YhZ
Ccs28EHuSqTvMNwNrzi02dI7And9B48KWJ8yn6z4cz2CLiJtauLhmMeEbfvUkEK59WT5gukJEqLT
m11okd992TueyAz7a3xwoS5WsAVAIcZWGAmenIDE2F25rnl6uDi9zRaagqi6H5JspzTvULZo5RzV
f6QUeJr5wiGeo2d7mObnubIK4kFuf1Ilzm1espYuzcatiUxqoeESesdhYMiz+l8ah35plo33ZqZI
lHHTr3zfQMynBETnY3nzr9nF/xvX4MaR1sip77hIbK0hCRjcljfXcvjxamj/iXejoZp78/8+Tzsh
0e/hAYJNzftiNkJWFxNZFIX7l05Q1loCySkNzNR1f5bMoF8VtJKIPOhSnJazRlvhu1qzro1rirT2
uI7ilu2n4EZwzmum98mbUJwZ7veDDnL/ZhBwVB0QYLT7WLlJzy2e5hMKmZhJKMs14nwxU3qIZxkl
nAe3wK1butznbm3Cje5BLgbfBiqbLFF3kxsYbbkzxojrkOURNVRsaGYQewUWxoE3EIBr6kjhvHPq
Ta7Z5Y8uzk3/nSKoGlYCs3Guom3xyKxio7c0vNWLlSXdNZOHq2FRADF7a9lmJhmdDjAAcv0TrT/s
IWQ/7aijU7lVncoHjBN6cziBDqNk3QKtmdabKNX0MOW2hgicdpjLx3iSoDe0GvQj2FhbzEUTINw7
TA8uB+jxRQWX0cY95FCUpRsWIAoYifWVVkT43qrTDsQChyVnePusPtd81kXbhpx4FiaOaRFmbXqn
6OUg2L+2GZHZq6K2HOI3mSPy50mXc+FoPUKY1zluvQpGXwj6XVcvp0nBcRnmpfQ0oY8F2u94cyaH
I2Y0gewW6i792SVMetkEYrRFBlve1wb6aXXfhIxevTbrb3SMXBrWiGhEVrzzeQFmwRPjSyTC3aqZ
4K/xEyqOqzhX1gTM2FLRzCH6/OvYzhVoM1f07+SvCSd/L6KHRb9Oqeq7RIvezOD5VONKAqqMIbTc
Lx1ServPHiQsETbELz2rZhYo/+elYxWLEgj/rhWKNOJStxU1uiHk+k4cw4QmEPkI+QDpt31WJ5yy
1PxguzwLyDkMTcishoQZTW8xIYskCuu4wdqJ3hYZnXTDXEVcskCFNSiTjbv43UVHhfhBg7sIXBqN
jgxqmanFWSAPWcaLzSQi5zCHGFw91ek1R8WF+kYOA2MxITYvmWJDnQu3xW2aJTOwYYof+Tv2SV0O
JbIynkN49DSCLqOjasapj/N8mNZoFfzGzE4s1EiZwtnM3rzYXgnj9djlWolOtGz8usEeRvYUyeFW
80E1DxVnge8dLylMt/m/ByxyMsLR6tBMRYI7Zf+R96hTjiUl6ihYLWvePn9PMmqomJyyjtHqyGO8
FUzqo/f2vxcbs2OFTQ5aQmm98VTQDkDk2Et0x3q9pohJG7U8ooRy3WBLTA+ty1TiaWpFvBKq+4Yx
k00nb7Q5itZOFz4oqpHqZ3UwLX1DwoFbkydx9qkdH6jrcM3qFHmVPDZ5mDzVoDMIgURvp/h2w1/L
nuADCatbxyguCSugusFNKRf/maWQwHDCuGJVws6JM6zVSIQhXUNXUC0v0EFtQHdX7vH7dtNMw63t
KCzug+YNGrzgz3bRi2UwzzRCRa4MgFygdy+YQGQGDhAok+bRvUGa10KBFWnN0upyF0iExh8kjXzP
D6s0kxA8E+Kc3jrVn6xL3M5Xc72ETs+HQNR37ZvvULHhINF1zKWLvSTBO1cX5yn82655POfh4lsa
Uet0mguNbxxHtseqg5Y1qkTJ4vVeQKpVz6vJnibvda5ubhcTJSXp0ZCI1gxbmSNj/n0XV00zTWI2
u+2RcWDJt89ASFnLe2kMttXSLEDb8maMFkifW0D1etRWSl6dLhJ789j0AQM8KD1jkIVh1YGZnofD
4tCyh/zqRlGJVwkcTIiEQkChYcapbWPQ5flvzTUMVUu1feOuS4SVBhhJrGtcPA65xT7OJSGqbEY7
hLV3NqpvD3wxbhvtWH3fVNqW6RfIITaAsA9tySjHc6hfpHbENkKywUohZJOTUjf7YOdb1M6QPcRr
10oF3Z3Ymnb+fG/nDJN9SqR4tt7A36q4BJfuO95gnJe13wk6tQ6gp4iAwnqgBa1eIzsNtbEbvBaZ
PIc6la5v8WHy+BUAXqiL5nyrvXEMWUaHz2hZzgingA94Pj6d02Bjnr/rme8EDPt2dDKMx4yRyCfj
TVvIXg4ZPLUl4Fn//YQEtBDK0+VK6aTDtt0bUq8sME2IGlo6+PDhvSTYXS4w8yqyWfRxmcOeInhw
1pA6Tjqr4nQUN8VOvbUuDvuo2A0ZZxph0twdvUtbkAs6WQ+2yJfTlfVrYvtIvSNxMx9laX2k7M2O
9MAxBGTl6tYS0ZCDRZa+lFYw8f+3BQZyvNfFk4xfa2vsTZm8QJcmrGZA2fAd4EQpUY5RDDZGrVnO
NB/SDhTQrNakug2b0WUnyf3hclj3Yg7HXxv+w7V1G/d1zGWyJmhM1pUGeyJr9+2BbRqiXvXDenO8
hN+PG6jX6a5XG9xnR627/Q4LQY2ntukeT+sR7NVHs4BLrrR01T2DLlYdXDogLJmLOewbRQ15gdrs
+IdWMBwK29JTCnL+GCYt3ZkIOncDRCfsKLEBSN6L47gyhC/s8IFHPy5J5BnuX6tVdu+r5MBigoe8
m5SzRpbriVySr/0o3CFVF5svbCjCfYCjRqjsRt9KOBZln2m84fxpnHBncO40+EsoVjyf/LKGq/66
xYcIHW72wvGiwKZ3QmPriiorhc23YW9yUWrnByt9l+caMFaBl9Bb4+2RgEVIzxZwT0AGfaONXXuv
VDIXXEYratZORNXVDs4ALSeWbNcLDup47kTaaT5mrqxC++6KqflYB/17j9xOZ4Weixqc6Kd2yyfs
y1CMGgrGaVaDj08DmbuqCYUkyPM6kFD6NSMjk7D97Lc7Xh+Z8YA2T6iWo5J0b7WVdBJq2Ygb4NYl
2fE0FDxSNAzNe3UstTpjZSBbRW1UPoIfyJyDtqSUiW5FvK/uYQXqq4tYv49eB4gfLP+uzNwQRFWr
Bpb2bE1ubjGo5meC1f9cP9PygLCasw8+ViA6etn//7teB24YQ8gGFYpC+4JheofPV3j3upkZ3HlL
M8OxUoJXrCR1cZX58bHfa33yuZxIEo88V7blxI1+S6zuL16DF8/kLFuWvzpuUBH0U2XTnOIo57UK
NEHT34o54sTBvMqzBf2cm2XJU5PAoB4nQcfIdBYTGi1sB8Il62VEp0AnjzcCZKwd4yAmcnam89dq
3TggHrdPlk2iG0N5wnqcVu4nF/+1Lp3S5/WRXz2xqZjW4n2Pvic/UC0gsJk7H5e+KrVmf+uEXPkS
JOZnZDHr/nv63FREzH9XQ94F70plphxUkuo4qKej470lXgfzvafsSwF7UgAebJUWt/HspuO7UX4Y
fy0bMzQnpI7UmrnjIAgjaNa5nSWBCnuaYHgoaBVWehbW+72yozvJ+rHUaeQ5cIu6ZZ2C4GI/42QI
k8z87Tdwi8HVEV3zEPrH4leQnoNYzBS1QNueuspKoZheAqQeFRD/RhoCygEVIiOhV+s5fw8dfud/
eSVb555BCix7pmzYAeRWgP8jYPV4Q9FNjCBsezG3/C/4tXC3xcXbNFEjVMh1GznocX5B1Z9lNuSP
pONdpYKgh5+VENnrtrWEio0lK6Uq7SI3fT8fOTCmYeLO/7QpPpAn6uchtmfJt3106c/RnHjxua+B
5tZt90IKwojxiLl5isrZ+SoCGveCqZtn/MhViXrvbxQ3jutpZLND1xrEsjkec3cz1FmWr7ZB/4wz
AT0goQR2qeqBnDozfkAjwzRNmq+HNfcXa03SoVZaRC3LsGk7KD9h4CnQU4qZ1jJYqa+RQDOAiCrh
DGjUHrhuiKxKtAgS6mEC1kdkdwXiGYierxfUjHuS7i7+0MqUFPcqE2DxE2/Z0qMDemFn9mZmfSWj
6LgyZD+/WfyMYRurALAb6GNn2UzBxmQpHO+a4spndLlDfNeUI1Kw6HjbfqZHuctH0dvCKQnLRvw3
2b22qMENM5A1SSy8DkqO2L17nPLB+vb6KC6KVZCAcjpDEnxjrcxChRRCV+l3HAexg/y3DhbAxKEG
LYFHWloEc8AepKr1w3rtUVwFNJ7px8LG8REJ6R4v5vKGR5VcJvV7YVUPloqp7rW1ugkIQ6VXgcf4
bhJR71y95QzS0c3e5dCh6HvGXP+YSU7wzsjBBFpNuvrV45bdxzgag0rAgc2NcALIOCDTGJl++z4t
iSBrS09BT5xi4KGqWbEyZsKGRAKiu2o8EKJb1Lrxp/LMeAeoONySbxkpW37Jk/PX9Pc/oSuggQit
mbwu1yn2rQ67g+I7B0mOaWBUy9rsljHUrx8VL0j/YRje/tpTwl1FlHtqD9nApMi0lThg9KXaWW0q
yXF+BDAaKvU0GzkWX7m9ctW+SKMc2H79KncPpZpdKBxfw7ZAq1TNRvvPy7WSQGITjh6QX00g3qHP
5wr/tB2YEr+bRWQw04BjqtN1kb1l/kFMIVMtutzYikOSvNzAe9Qoa2I7XNN2pwTAcMy5pwGqVq29
E+eb1MyvSUDbOPl1llZFPyrTJr2zkz+pHnjPVOssbDkqLbWFS6JG1VJ4MgNYHGyN0URRhVrPbejK
7wIrv1vi6fxTviOk+PT9v46pRraP2aMj8wpbz9esdoDt0rm1ZFMwurjFMsp3A1C0unt9I49vASxN
NrQWbec4V0QBtjLfSC0vXqYIoZXWawNx7UQ3EcGNm3z4ej2yEcE5sDlvaB5C9EoKq5I5w8CKZGle
6z3+obXmi3erogMCLjTyrACoTr9vmFWUQi9oTd2GOfcfcUe7w/mStj0pfqrG06eaWsD15BNo9QXW
c6iIul86simMJoJEIrAeeTj0GeiaqTUA3yEjlJajIrWpGh2Fz0ISEr+okjOM/xmQz+HlUE/Ux7qs
eSrph7QCt5MOFOJyMbp6w0QWB7NfdzFlokspQzoliQVxedxyBQbdB0LTLruzVMfLRWzr1ARBHPTr
XOXETrqqYVDPbbQHYPRZM/Hdbj1LWguzM7vVHg0zafshgixGUkSXH6kHRVIM0SxpVb9XMpMX27XZ
T34PJWxCEVm2IHkb+kk7PS1eN0vcbwRguvSS5KxwPzXtVYkV0dMCBAaPu2r+6FW0IMjMsfiNwdwk
cn0wZijmZOBZx2+Xv+I5dPr1o39ps+7A0DTj4EssDBW2szWoHN7RM9luNfcSYrrR2q/OGU30Pzhj
nChzCqu0Fa7Ac7vOCjkldLhhUu77Z5bwolx/VQ6w5fj7gBYXMgkK3oluji2lwbEYimzLXkfx41y+
HO4SsEAShe870U6OwNHcmQHblybtLPMsPANBalkwJg0j7rV3LIhSgP439d8pJgOjm1oFjYHrKhCC
Lrs9awTB75Hz146v9NqsqUBVMBEiLQpdcXiFhLSFnCJr9KmW+bbKir6zR78bnTNFgsME34i01uwP
2ReT9z37gcDukXt3w5O5tYiNvOpMzBMgm73dvSl4u0Io2ZABVY/B7ChWI6mWhpe0w8eVRrA8XWce
BZilhkVCXsvlcQpk8kw3w+vCl7c0Hc6+Q594IUfOojpsG1NNA0pxwIAC/rCll+Ha3NApqAJaBxZs
Qhj57sU+8uaQjtf8CzGsDoDH30MeWT5PZBjOD5Ig8vz5EFJHtmE+lgAJxwm9gKNepw3wTPke5dgW
R99wThe1x3JsuA8DgKfewXCwTgm4xG08vyD6703SXQNg2z9/kSW5XKH2ZkcNZfHA/EXpaCtLMtxJ
DjnWfeYt/0yRvYDkv5X9qMVIkElGXDPafUE1mr1Me71o3B+oBOwmj9BLf9YGScAvVbyU5zb/Npwn
lJyKd+Qkj6YCiAAg9D1Xj6EhZtTaTp86Ki7wrx4Wl1vsMryAtHFXIlld3lY7F8KJzAOIFMdn7P2P
wEpqE/1BoqWw0iRLgbjBe2Chco0KnPv+tebugqbVk3tty70iEmEo7hdxPe/m9ncb//aJilqQjcE1
tYWuFIzS49QyxviumYMUtaSGKXpEEmh+tAHQ2U34Iv65Wz5jwzCqOwjtH/kxZEN2q5OqtcW6wwhE
loJJw+xMGmn2HesWKE924chALIdKqUMTUQgzF+zCQPB0BXPnTlHy77GxDS5wKHfaM3AdSOOPv8+x
DUCJNS6CV8SnLOyTJNwv5Eep5RNqO0TfFtlQBtf+NEDN7mbq7/kgq9qJSML1TaFRj2b+ihaZ2F/T
kTwYKvN+nRQqlqlye5/qZMgtoKak6Kxxm4mp3VKIvl33engIydZAQFAAKYRwQJDb3gaBXYeVxkDU
GxNidGBmiFitm4tUsicvk7GiKSYXZqknW/xMcweF12NM/bKigbETjsIOBV8kxczZ4iAtmTAAZ2X8
7tJ8osILjqtYDe4+fIzmAzH9HWsQiTIHsDjTW+EAEApfvU6hGdeoG7DIGe1HjCJNs9GbAMiekuW0
mPVs36fC4YYUcFgpgAI/LhCYmDkisNNN/ReW3BKVTScgo2ksUKOxzY7SFD23VeH/7svLkPg0rgfT
u9BScMXRUfCeoP9HyGIKQGLnTWGDGs3k4B4PZf1qnurFIIDwqKZbXfGXktP72ZueL9cNBJj5+2b9
ogMJd09wb55B0TWIu91LTF0PXY2APGGBmCXUA8TppdXpLKYoMLEtMYcHjg2f2MOXxrX93o0J38mz
YoSfy/02Ij+93jsEKrIYdc2Iq8Fwxb7YhTilLXoL5BI3K+6qhhs8eWZctIw1NwlAbYaX7GW8lBKA
mzbTXJmsmoqCIw8Fcx46YTVVyyVZY3IiW7/wA2nVSfg3yyB1I4FMsW3nX/sAF/d92D4Q0wfkapFo
IqIoX7gycHbYzYLZN3U17MUrRNA03ABGKkBz85sYvPwWAt1qPdiYvzZKex+okMcK3dK0tPR0pGZF
QzQZw0iyxp4n+OrfoI+tRAxFsgkcl22XKrn4L+uRTSX64nwGbj+R2DNlPSm7ENWDR4SvD9GkAu7V
0OhjWFR/Vd92YK4Z38iDOwwk8noCdo/LbwcWr9aF5QTb+aqnuCT8ju9JZHFn+1wuvcOly7yCFX7L
pxbGjUc94lrVKeNdmCI6QYTMG7KQcqg1g8qbRXccKvmhlJ+fbALvwWWnNsDqpHdstd3GnND/MWz+
RMxDkmQW3XTuYmZW9mdsF4m41rdjW9jhgqftPfOpFj2qjCKSqIo8vvssKfM7zv8zVa+Jyhmo7TJD
QOonxeaezm6WeokSGctjTU/yJCfxijHjNN6HUbJPFuHVLWN+WjPcJ8jTm9TtNUpzq7R3WbzsYL3E
M2D9AqaySRX383G7S6oPBO79ZhnT2iCGi+OlcUdgIJ4vLIPG6MdgXaXn17V3GsfVNilZHZ5kdZHu
k1F4CbS/XJGR0j8C5pNvbt7neTRPYdHfkK1jue2w5iPSk5SZdVwet0GISctyWRgB00/y7AWapFS/
49RTska9igBZXo3Rv/LLzk6uBwzIFA9NzFRnLF6MOqKAiMDVz2swebzOhCDzJNI7sxO6grYR43Zz
1kPt10jbTcsTrZluBjbHn1TaKIP77AquLX/faySaZoVdhcWjww2yTib7V1OXWPWGA/9heZXFx62k
x0qDaQ5wVWwGqi80UnQGy0FGCbek6LuWi1OYNEDFb0Epkl1BsZ4svGpSrV5FXvfVUUdk7Y6Wd4mG
CQFWkh8cSXUsHdqcX0S9lpJ3vA8KF4hQcQXglTJbgYRsBruGMcVftFSwkN1LuDkh20w19BYkh2mj
5XG4/OAf8PZ70Bs2Dt4Lp2yX7kKd/eCx6zIxAi7K5DvYxMPxbD37pfL0Q2FCoDAFuj+RGZVcdYEp
JSjcAz+30DcK2LrnnxYMajDxQBRHG1okxmeGBleBwfPnoRXneFFr7/ERZyNm9+8E2J3ZfZI7BYJX
MdZZKh3Lv8WFHq8XwOTYBRguRNp76x2qBQd6QNYwOgqe4fI0VIV9b7Oehd7OIY33x8HuTeeYfnea
JxIiWJbigIS5290Qsedb1ztj2MjAgpqhhCPLlszxByJqO9a+oqq12998PfRracibK+U54MJxmrKk
I/Vmlk/LNVREVgzlLwG4Urk2FIFD/+x/LVL2EXT4SuJlL3swD/hwTmH6TwEXVvBewJ3iclzBSSF1
r6XVdlNySzR0XD+kDE8GQYxlu3NuFcQaY5CD6gkjxUPutVqSUTn4JDJnvpReEa5e0Bhz+WYLijrt
YkXmZ7iHv/LFmdoLkd1oAvBgBzzCcep8O9+F0jAEqi4j04CmObl/4zIM4VweO0qqZNdYtMhnM/MI
Eis+x8UYPu+3VnGr4q0fS3oENPIaXdSVc+nNG08Q5OUPwYPJjqgx70qsabsYOI5a/NXDjN9ba6mC
UWRrt/tES1sjnjfGwfXz2FJEIVuRKD0mdrOrKkWeG/4k3m8Or44tA8qRsleDB+ym1lXFeTxIvT3a
bndN5FR+XcH9fXmWmM+KCDKo5woBsMuprlg2Prsiwt8gUdeMXu4vBQUXZOBezGSyV7SP8DgMN/1t
0zsUxz1Glo9X+lFS49CM2tKEBBu3U7pF7AN3YgY5dU7w4xDfH5BNqLjxkwX8YTLd3ldZoyeV32I9
y9X/+VgL8lXGqS6Cm6QV5tPHiydbX3iDB5y9p/N7r/x+S9/o8U4OrBeNaWsRTyLY2c9QcuMdWRVM
NbNMjXGZQCUJoJDYWQ/D0jhEEnDwNXDWex43FcRmG+lKAOo/G+08dH1EgoSavKLJN3gz/fUdac/R
Epv6/K1d5kSsalHUSH6jXYJkP1VObH0DcHh9JxA5BVU9UfFyoFm9zkJq526zHlP9WzIJYaJYPllA
OzypljAu47+hiVIJ1z60fctGQfR7qzWi1kIbbrzZUuoEfSrWQWlP7CFHAVX5FG/k5lEKdn6R7HgE
hWTdWTMmAMZ2mpL4d+EQ/MVETXH4fGkAE3ZCeYuR5xMbI0LrkSFa/AWA0JebisbrsEAa2POLmyGI
wp1BhXpaEu3sOmq/qQ3aoAYZMqlccwGeMsZ2vuCo9iuBGyV3qfaNR1pYfZpzksajLFxPqXuqp6aE
0yUAN7+yHrKFCc00iD2s75W95VUy7gwLrAEpQekvyRgnhRnHMSFkt+PuhFLuQ8psmRCE/qC2ZQ4L
k0bJOYfdzE50EJNQtZm9JqN3+X6bFKmpRcinO8kPlupBHkPvAS1Ax/9ulCaJvlc0VV5m3ZqKXlA2
77IbiEA4i7Py4wuRzuqNaHqry5qHrysu1PG1csmeOCZfqOOzecvJr+MbM8N8Vr6tZE28YG3G3aHR
uinpqbz+28V07pOKK8W1jrhiXqT2NcTJpaFe5hmBmnYlUX1sYkfeHBDykanDOAC7hGmQW/VW15kJ
KYaMhjP/M55lsHQQe7pmDcCworgRKKHdtQgDDT/R2J0TrMsyOZbUfma6xzBoLjq3xyUb3JB4vg0B
CE5hOI8TEx015HxkaOMiEquUYx7P7UEzy6BxZBPYkbXCeJSInEuDDY51cTfV2hDfwO+XUsGwp6ru
uYMuvcXLGrc18jVYtFDPe5I4luK90NLgRMflZiKwWjHK3Y+pDUnN5JkvPKzYkvUnOcaTC/hPkwTL
+m1w7QDMxJc3YI4d3lltFuKXeKmtNhJ4KIEpHT8Ar50tPq7H+a2SlzPvVMnu6cFeOklBu+OVcwEE
a6rL+4EXEs5HrG2LiXRTDAOpToE/OaAGOi1XvInudgVknUrESosVHMOrUFajmQiVGVSdXPw8lzRG
WT31MjY1QMkg+rwr5HmUBg647Lje9yl9nVtqT+wtRfBjNPtg/be0vsgytLIvjxY29E9rZDtjFcYn
8qmpLrxrjOl77dcuJVqjnep5UYo00JbuPonePY7NDW/K8nSwxQRI8xhmPuEKLgdi1yurVIowkc2W
eoyctH2bRFUaIr0juOJe2GdgTi76Ap4BCIPese3YADiMzM4a3aK/+RQbaRl9IiNj1shCk+TSUyr7
z/SdFtHryrnIpCX/c5vKZY8UNAmddLm9DhBWOTDGWMAVW39rgeZFlZurTqvDXRnHKdgyubP4Ka4K
eu84JV0QmWW04GFAWlplik39trTVb2ooYPnI09P6ehC18Fa+nI23uiszymc5MmTrRn/v7BzMcU42
BLBt3ue3Ez0vmV4XLgRGMqhxvrvXrtKNTtFfSVS9DD59bylBkb26H8ARpxnKnkBAk5ec4+LfCm7y
3ACwatCZKfUYZHDSyzqkCfz7ctBEYmPD34RkyWAiuaEmR/3EvoA42LwvP5iKrZTZB/yvfglguXsl
wbMzlQ8xAR5Z7I9auLbff8uZyLTu0xmkGhzQDQ3SIgBtAQWddtCfiqOkZFkm/pp2bk0nJHItMKNH
DujcrWpAU6TnnfaPX0vKRoPlrC5z7yUoUQw1SQql5rdIHJs+cN2OmnKSfiLEe3m/Nvd4y+X3ExuR
31kF+pqVDywCBKETdhYsnt3GOx0bU4vit02MGcBwz2hciP6r+c6U5ULdo0NdUIv+K9xPxsg0+vgs
sfI+kSO8wmks8T4wcYyWebxDa2G/6/e/Cidb7OFOF9k3awVEYMVVCIhRfLdQriie1oJTsAVXBCzr
Tut67csnlBeSYyq8pleCzByz+wNy/Q+8ojVP00FsCxHT9j/ZVHF/bMkYMy1YYxd0+Au4zRQ8Q76l
EiRSz9pSDOC+/OEuBdXdg4suBqAVMsjflAOVzRShhCLPBvsMi1V/RUengWI8bNkehWN+qI1v+y37
pR6RYYMK5fsgKNzJcLbtQe17phmk44N9iZNp+Vuf+rJREkKdu+NYIdBlbO78duj8vFWalBlPbEuf
Q7e6Wbio4cSvpDGaVykRdYfUjBw5/hEaY88y00SIojxe9v0z+in2mpCkRzEOAGSP3jASDbRUNJv0
kMiG8ZiDvVJ7Z49FfOmASDsn8InpAHiMeTr6i4/mH4OW5zqSY4Tm4h4aAqO4k8FwfW3+RvjlcEbt
EI51fCCEub9IfVltYXZv0jHW2xmbkYaSoZ9EA4qelciXRR/UtP66nYTP+hQkZ6O/+5aFSQRHYOuO
gnBcfkGQ5sYra6irTuY5paiLFaEM7nSc6FIwoSP838llKl64yWZSWXAalimvPzYkxhWCk4/pxp+U
2N0X+mgqTJnGJIytnc4LZmAttke513dxk3NK8ZHvZQJmzm2k6aYOrGkQ3JNjqp0a863WZ+ZG5buI
/iV3RUSFHI1tYMsrZage9JFu5siX0AdgmD2nBq2+vn5g+YrlETsjvw6CI/vENegmHO8ZUnWdjt1P
sbdOp3TCRZFaXBu2YawiXfLW98L+8taLgyKTGGtx78wsuS4cEqHGVLEqP38Tnc88FofTq+lyj04k
szynHu8O/Qzc+xxih6I65Qh4flhn0B3Z/ikmvtmbdU77occDs4RwM0vwg+5RZ/Jq/oHfIi2kD9gi
ix5BBGHAVjyfRSK7n3+HP4S5Iayubl2CFc4rw1yr+9QWtppdvffrzwnYrnXpiGtgdlfWVRBvOuVY
pOXW2dR1xC4fb/VBV/rlKSJalFzuzrkpbqKWiJMtumxCTzRb58t3A/7H3xif/Xf0Uyz4wkA3kxDf
s0TmSM9XvUaVj7oOIa0HeihKn0Gp4179ClnsFZOaR+40INE30hpoQodTBt/3eCvyCykHG/49XrQb
YWw8fTS7JdxESVvq20NcUvjfpIl7cJwbKvEb05LrlVw+WJSq61jlqSGRyYUITzO1dJLDqMijL2Ju
xHYv+HqRj/t4fnHx/1hp2pfPu5beSy7p3mlx8XnhsO/LhemAVacrSBdjbP4n5id6nB6BZezqOfgz
yyhd6Sqz9K2fkk0FeFFXeE/fif2cxZElElPeFUF6Jyc46akwBF2kZPjsGVXFSx0yyQc7Klcag1TA
JU03kpREGUJEyNwGfTftxrTVhD6GCliqYe7f3vHipXChX6IepqF+RQ1OC334TixQy2VFmnWMA7BA
7rZ5Y9sGxvLD5bGHEianrHVbgXH6d1yP/DzAWn7EYxNZ/rrgm5kpvuAxOI3GQfR7g0UFB8lM0hAE
lhVDBZz/A0rV7CAH6oS7v3bUFbExOeAS4lsifAvcPw9YUhb3RjWYRJWxJN8lShtBG8oD2aiTDGro
n70liO7AjbM6oGJ/yBendKcu5BWu8XSxE/nF1Zj+cmz793LS+PzCpbQ8XKMF9uDtUla6d6/kasV2
6kihLtDgXlfw96OErlnJwtZn11y1pJaDrxFE8mM+I3HqzsGq867K+sVOgbS4apCvKdAJPXUHG633
Pdi4Zp/ugdD9W7Sm6xax2GAwVUoFApbER08IRwV3U3wFAdcpZqw5GU7AMVuQ9opw8YKG7JIY33RY
Or3tbLakL/+MG0gj7YoBOiaKXjE+NCX+GCQTsW/dTs2mazDZ3txra7LU0xFxQ+q1oRmsaqiz6OGH
BrZkT49u6kJ9c4N0kwShFewKVF4ppyYBgDkmLjSCXn2CpZ75E4Wcj8tN0jKPws4ikxVH303fW8yx
i4pcg4lUzOqjba9BTlSBlALmxWogcbJCChzXDY2CFgvMKgQhbZuzzkb9Rb8lbCe9Dw3egV8YcjDM
RedYzM4Bnfdf9PPKwp8cL44sriUImBE/sMCuVqyfHK6QHOQ+j9Y2i+ACoSGhx/a/p9f7a93W6Dh2
32j1Uno/L9/bJ1E/9BlXGsPiyBTIgAKKcwsI4S95LI6aXMPfmAhTXDisMRrG2E1bBavzMbJfA8pS
VJBkgsNPtne1Y93JS++8EWCejAkXkGHobrmjh1uVbr+BBhZOcpnXN4+LKCi4VMmeARkmjetTJiqn
ob5eS7bwdU9Oj/UBmu60iR1kelqzk/NZTqzDFEWhDBM+O6aStb17h2dldTaTVvZnuNhTdTH4v49t
9XwnfjzWo0H9ooBvOXLJofrel+jt7LzZ39wk9YZmTtkOljdztXIYZHWa9Y54PaDXs+Ibc2RY+db5
edllcBh4Es5eyuIqHC8AIS1/k/ojLd5Q2HMQM4hqjHMMpDOZnNMs/D27nC6y8FZZ2iuQkh+nIfF9
WWoRFLldR/9nsthGtIQj7s9T7siW6xi7+QL/si4TkHO+H1LWBczdvTHXhCh0aoZIAcmv4ekZt6NI
JFO8EQnl9SKb51AGByTyKQkoexRRMY/aLP51v+jaKUknLcO8D3FZaU/wgmmszxjfyO8ZW0J0C7pf
UwN6o1mskTT0Hzg6S8yXKxNPCe/Qa/eKWro4QNWPr5DBl40JWIVMGepeJHIESvjlQVWcdTtmztsV
hXqa5xm2CAN1GAGAiKqcXPQ+SohN82lXIrusR0rQVA7opgH1Cvz4VybEHy7HezdoMqA8xOUZOu97
2/wJy6Ier9x8X6s88Apu80D/ElcsqG8sjVgD0FeC8F3d18wRtoNwVvVYDk11NO6jkPFaCLbZfwFU
ptVpHu+JeYSQfCkSnzd8Hx2xjalyRkKVvHzTu1oPasfKHS18lATG9M6+062jh3ImuL7nA/S2s7mH
oV9MpsPHyN0FYlPEFzbOSzFN6+6wPCxUW4ktu/gf04iqcT3dFnUkcYhPuC991TzcBHzs/DL4Kwsj
BxmiUCnJoZkYpcSXUTbryqCO5pHr7gjMYDammRii3tr6nANn2TFsmyXPPm8JNMe8XuKHVJ4ZHdv9
3ByE6Os0LAThjaGZfbomCAMgqtSnHSm27B7GKuDW0TmR20xfZjZRhirCVBWig3/dfkY6NOFsybw7
93v1Xqe6PQene6J9rBpYZ0qKp44Ft/VqiH07gZxmfeoPtOdld3JSvWpNKFK1STGrdAnZnhB+tazZ
sY22ehu92RByueMVt0RoRIl0ll755CDqcBamlBDmTnfZrb1KG9kDvNHAY6vwADJSu51FJSHGyj7n
2mN307b/DdkGieZtF2CTrYnDeCETuweekg4Vb/PcazTUMEjfDFVTDA+BZe4jQGDvWuYi/M56WQfu
FHxk4iWl4E2XtYrNRFjRr3/QGBURVotSSG+Yl/tBce8eeLxG3gVbCuRDpngLDRf6j9znApLH2Jd4
97T8vI+FqU5ng+8Uon9zhs5b7AwXE88CCACGXSqIdJb1LV4KoEU1A3+BKmI/fIU94RATZ/z839BQ
PrdSQ3g1EJfQowfFAMLIjK5Pjk4P31yXDVRQpRrXGO0ZigpM1lz+J3uVbFPGBwC16Q05+kl6rR5s
c07XxtTWxmSHNqnXVmXaLizL8jhdjts5tDbPECoKl+ik7Ec7yMVOIy6RV+PC8+SsZJlrFY5S2WJ8
kqu1Jl3u1xQQxEYAbFr8j0xExCVzI1yHuNAOhDWBPpV/jXJcIc4iXgoRpbc/s4CIcmaJol7zqnsV
oDOTSX440C8QMqXrUjRJ5OHNyGuPL3N8ydu8ceXnuKVUhYJdBO+pLKBpgs1SWO2KSsk6pAJ70pLi
rfgwfkz9IhMvqDyfHmUnNZNNinGCzx6zXoPQEpxd5+Ihh3VwuyAP++fl4/S4LrAu+PWiXYeSPcpr
FAtlfIAIpdfn/EJM0HuT1knkOoZQE2UuokharZynH/NW640apuFUai2TLsD6yyQv9uqy2WfbLDPd
UZsbek6DmNj6BuINo9Dnp/ef7dOJ4IUk4lf9vffmAsCbadm0Gys2M6eL/9IP0XPEbeNMvXi0cJ2p
t4uWrUjRhOKfV8ceK+IGzIxrfFai6lDHWxEk8n0symT1z7H8JcHxjwndICG7j0XWKK+henUx0C/F
xFn22iBZgkDqF9sWtkjzsfsv/uyH7de0EVLrHL/qCAq0jOOxgvDAk3jPHZwBBhAdMyfd96qRcsxv
cGKOh4E+sTBbCshrJY24QC02RahED1zG0djtp1smWoTp58SeY0b/UaglMqlzwF+1yHa2qfIBzkaB
vU8mbKTvUB4qeZCAUldyZxA4Q+hcBASM9AclS7NSQaRvLTb+ttzUi+MbhGDo8r8X2YEzsqzVIPZh
GYiOae8jKXXxLNOzTlp5HIuwMW0zEjGmLVARUM3nC6DvpvBXVXfex1PabP63YXxemG0EHFX8WvRb
SjGHEeqUj1kanI+COKLnI2+VCna67CtS4xLGQYUQP5/Ux2ldy6ly582r/Gvf0lkVNfFzDeh2zfn5
QmQpw5t57UxzKwmTRROKT690CSk2ZVd3HnYkDA2c6QlDS3PJLVi+EeopLXA2/obWGsiI3HDaCc9h
cMnQiyPgnTr+4WTAmJBzpVZ3E3lBljmf9iW4STzGfdQxZknV/BupstWZHZXjwkXNdjzo35yY08xO
48JxhZUQRlyh+VuL+0akhaOTeOt/TUwJUNbq7RWoFBGGMLimd4uWNeMSmehkmExlljSekamkXlqi
pbgFkbIpGR/zkPvcVSicYCG3RE3U7hllWQzoTh8gMiVcjutL0DEgZxAZbjmsjwWClbZ1wYl4floX
SL+YiIvNQAOfw0zI6po1Na6YCMpmZo2k/CDimqHRoWMYHLlAsWrCcFhAcJ1imhwP/zyYAPlfIGHm
emI+a5OTyLP11ak/169XvXZzbHh+0NuNnSmSpyTMiWFh8T7ATuBPfVhzw5XTuSUZRdsk7tjpHXW2
ut2snw7dlFWHKsEfYOKlkbrOg45+58dlG4ypaac2h4D8VKcmTIDp7A/mvsaqG8N74q4h26yh+9p1
jwk+KYdfl9mi6+ftreoQ3ujnB/rfI3/80INjy7IAAaFMHtJsUArr6XmiFrzRquS46d7NbwxAEqch
5u3i8pD+XXAAh36Zqa1iUo5I3dColiK25OBiMuUEipnkj1Rd+Sn69wtH5eTP45zGmZzoWiEhVC0o
RXO3SoZ5aRQcqCbqU/C621qJcsQ8IJqpigXbem3DsIeepDGQSgMfki3xuh9prQOB3dnegZLme81F
9AVV3jrxmHHbwmxkOhyUa/wR6Nz4NTylWwl3kBFCVDAHfUzH+ojE7IhIGPiuWOf0wo9lLvc66j+I
woRWqOVM/jr5bgCrzI90IudAz5XJ9mcgbuYQerST+i7QfOlsns5xyy9Fli1KRT0u7IYC7CeJUOlR
nryehnnoXC+gZgES6N/Q5AF2kEj90x3jgKZvAr6N20QqIRhfxGQSD0O8pIfWR6td7eBCpMBroMOO
yQ2CAim6PUWOiuwzVM3jLBxPc4kdnFMRV7D2OVP+8PfSEy4ID/w2HEsQJP1dvCgKuGTgkDBOvuz7
Ag+NRn5SOXPwrtCYYwTRMxuuviLVRh3cvLFgFcPXFDAII/wZandt1t+IFE2GzbONTaQ73G2/zqsP
rCB8aBSfjHeQuvix6vP0l8ELxouHa5pPBzSCvo+TifotqPl0YKMa9baHdPL9nwp6q63JYHPClteI
Ie2epRA0VJ10cJt4hajCrOpCpX5NQA2k7b8wTtkmqcdwgOk/BU+31VGzt3Vewacl9kxC4uuoJBbl
u4IJhT93bd893IotkFiRUskUl1l6yukM6IjAHayrahDkBTKZvOSDv0CmBs6hvhaD+V2HaKeWliy9
JdusBx0dH2WnlNBAPPM/Rw68SzJzgTLZYaUll1TKbfxQ3CfZDU+F8/GMLwqBDzoVjFsdJ800r96M
R/dxnfuAt1Okcu7k1gfcTZGWOLEHOr/5cR4jTgBT/l+3dVoND5ECPMGLarb0Fmy1VwbBlMkFgfC5
T2ZH9WshsJA/d+T4gi3SYomHoIiuxov97wghiOtc3p70n8mkjBteJ9552f9mBPws1EjKdwSA9C2c
bkHNtq/Xj6aNH1qGj/8BTHAbmZewN1Dv6AlIVsq7E5Y08omzBy6Wsg32sW1gxr1ykWH+yhXNJxz1
DhJNBfTZYGcmdBGvAjpYIQmJRJ8iWHcCbDUD+TLkeRQuRAMosHRAuNBoTW1G6Qui1UQGctf4emlj
1NTCIO5WNGan8pIsa4CJUqLM+tLFvQNjCXEjpJnxrRY0f0NIuMNfACIf+gnpHzhEokiTf8XSjHZo
anspMWaZAaYeARTFJ9LvtC7VI49Kcro233IllOCZxDKvFr3v3FqduRxtQjcHU0WGtbE00nz68F+v
1qDAqJQTQv1S+ZR7/FU9eGLzmubZqHU7qWNWE4RNqBL/CnUWUjDc/LtyE+LHAZox8QBk/8wiIpEr
1YzytBIUvAxweBnaI57z1CxnTi2rnn9zliPYOjqCoWJY+syixVOwWrjcs8nruVQe4UXjeu/ICVz+
18CaCl4V2E5TGJo6f2ENpJt+X/KxYICMLC4P7Tv1RSrILIRWp5l7QYtGU2/uVUaq7FGPnuYJGR/u
r8T7N40etNMVfpKuDnhr8YG5G3aWCiBfyCN7sicZ0ZH/I7rAxhBbpjGkN0lpDAPqYh1wXDaXs1pR
L8Kvn7ygiN6L9ckH6CR1HQHB9RsHjXYDQGp8Fa1aQTRC/+IyAB45BBN5Ai4u7F7/mebukuItk2tO
B1AFSUGnoepfQcZbAUuqL80Q++CBnbUGhwsqx9Jf4OOjgl3KjiFyNrwEH6S5SE7m8ATVeTu2OEFg
Ch6PQD3FDpPhuKeW+9LmSbylXlUM429XD8WT9C2EjO+P/TT4h+zXNdQq2k5L71MtMcQjjmxjgIhd
v57dhveypEmWmBWGVgPzxgRzz8i2Oc20sdbmzBmfi68vIx19wAYGsGkroT2tml0CFPQeXrBRLIYa
9znCS1bD8SJC3rKwDNDaQnYyC8sCrsTheNtaEB77oHAU2g2c3/1FYP3CI/BDebx1R0qZlIkleuiP
KKkWvAyEuNQdzLrJOKKtJrQQD5dcXm+Bfra/VTMeO7o2AD5+LJBw17VjNrAn1Ntmv82HTi3+Oh4+
rReALf7j+AZRrJsb1X7WgJ8pHRZKSnnLwMYZTAWxxlacs9q+8c6PocItI/urpW+PHr1aVZxZJpZf
DYplv43Sv1Ue2knE433eYIx785NX6L3XrMy5I4HE23zjbGb62HfHPsSKa+rQl7sXKRKSsRBLJq0D
MxiDVsh75fS1xFTRicb/Z3g2C2n5TxTDvpRvCUkXEtlECb6my6BgDVHSmTqxg6Y06TqjLYcgN9jr
95VrNaRZ65vcgryeE06FPGVGlp6O0fJIQ/8s4Hm09lruvad/9f3r3PbxITro7O3AyfC7wqzA2Aqu
WCVzIlx6JW1ii85husHMSgCVp2fquLPzy7wBX8a5rdMqbIdaa+53tH32wuEyN3jIN5ojqgJfVqkW
ATetktOnTG3vFOQOeDg7vQ/ZqlTiDLS9DWijv8o10KRqXX7j6AiXXTvB9eb9gCBeQs002vpHd+62
OABYahYt8VSbrVAU9Qyk7j6+z+7VhDEUYe5dUnkRYjEdU3VFEwE0SEaINdXVMtzeTif3MkFZRhcj
V8qTBce+pBuAtyXBhK5dvWARWpSBOTiQ8xpycOUCR4qaDCjGButHr807aRh5Z/UVY+EBS0CQEXap
rYXUkrluSJ5+8/clVDC0yo4Gb0nOrFb5ctGiy/PPWvV65XZNmOaFBG8rwlSTG36neuwOm/J0e62M
Z2AXrHQLrFwa/SjN/HLOLL6kM90Tn3wq6O/ZtkMS7JFNczBARJogRVn/t8Qpp9dsOTj+6iusbYlS
Nq4mkJ0ksolr6KKYJaoBhIgPaZYrMhwh/87HpZDaxt1j9xx57dggbNoCnb1OE7lYIYZSqlZELuhL
7ineGpQ86iV4aVQ4A+L+wS4tKRGUFajJg0gDXIkGWALHyUoHjncoaxg5jXl89cQJcS7FQXV6hy7+
zWlfOFHRCPK2LX7FTPp5JZdvVbQgrOR39fWWVpf1N3inKtK3iozqTxDTM026xquX7eoYO8vCxBm1
2gWRPcSl2v5YN4TqV+hnvfgmdCZFDDJ86uUCO7pepIQlNtBaR3xM9XjK552drAvloRI1reGaiX1N
SIv6gsicCWer8gXvOoafoQcN2w7/yaCtN8M4cR2mUFkmua0aVkc9VYkZmviKuCUXSkIYzg/9cbdv
Z6QKn3203g1Y9NjCO8IESQf14dYMOeAWyNRGlyQRi3StBov0vHLn1iP/qMges23Br5i0ziBy7Ha2
UunR6cYeDfJALfiv4QsTfDUTh+QdY2IbJ6h/1ngoWtxCUO4g0ZPnSZXNNdQhbf3X7ZHZOF7pzXZ9
o9UypmbRDNqO6rdxGx72B6g/9VOAlvRMCNaAZA+1iPGnaUEJ4bHjVwD0p4ejzuJWPfQsfdJ4llkZ
X6l9YIxZ3h1h38omis6EMyu8RQHPBxx3y5Mc0p35SfiqzsqzdhMdLcCbCqvbdn/6telDxjsK8ALp
bXVf5lORL3KeBpkJLKGQz5o9CMX0Q2pjbLM0bYEajiT3CCK6D2Lgs9czf7Q9aIC6qdD9Y6dxPJ1Y
nl9bPGgjsXRR4Axr5auTKiAIux/Nf8251Qd28+TC+CzRBLuFA3hjNkXQIhrjTXYF15iz5cKI074y
aDCPT+FMq5fM+UH47EQRL4211TLxzjFPVQ7YzvfWjeJnTW8PswCMDAIusExeUnZHqPv9LmNmIWD4
UFfp0eYCLQrXeAwulfQaJxX+EnxTSF1PoiJAN6VPmj4OufhqbFVGfQHhqEq9qDPxVeDAXS+VVxi2
3yjA6nyPI/6M6s2Bf0PD+ZXGG/tu7NcDP4lcLZxY3QB+Kzf4tf+tjPo5luIC9Zm7GdQJp4jP9aYc
Aaz0Pd7F4VNERpcEyBCly6FbwXOY65BrfbOsH79RSuu9oR9UeQy53SMxxr9pTr8PwHgwgzhLWAg5
2+zrn8BodXCpPPCcwxMrWwRqa4u4dum/uY/vgI2TwhoKhwEInkCzOTOdcwX5K4BHpyANq3vV76Xk
i/VhmJE4T3JyhdGHbhDyUjXeBzWrLHGGLzqrxDQ1ZE31V5u+xNDmbtu5i3uK8rvsVcSP2pQlRzsp
5b/aQ0jKNO7bd7WAqVVpCqIuprjcVvGV6UJZR2f0SiiDF9jryUqe3ZHZHQ428dXu6BO1rJmfamXI
b/NTjn+wqndP4F6MGiK9I879LxgIx1PK4aNXYduZetQXg2uirt/TwX6p0/tTh+EhAhT4nzi7R/MX
xeXaLrPQszL1Hd311q9vWz1c8gDc5HbnYtUQhfMeOysQpEOpfGtqKsL0+DJtCqBGxgd6Oqo/UBpY
mc0dl/DXxtQrAEMRKv05Z3nIno+DMzeOJE4viDHpxccObP/aHLge/PKw5MoCo3NE945/JVStrEkv
gXfxNL9k2isODdMxgBRMqWgs6B0P432FzXXt0jre2PxiKiCKyKvupVPkWDUN2FSn3oJmlYuGRXd0
cmHECdtbXjAEfYF8BNQlAveO1smXtMP6Inuk+wXlzvIRNbO/O0mdUSSrZn5/eu2sPmsX5F23i7tN
HBP52fzf2kel9C8rHjL4ztu4M26pBJLSeR9c7h36B6NWUkoEPj6nXCDPTuoKH5tIws9WH9lJ/RHH
yoHUbcCWPmX/FT4IplhhmU4Six49eyj4EFZRZsJWlX5QeyT6EzA+bQTJdIyl2deNcWVdPBXgZDyg
mhxgqScNNlAWid8YPbDAFaUzhZhcPXk08M5ZScn5RHPXivnlLkATiTt87CDgWRgENb2lfPytxlo6
DEkS2iwGgmhjT4t8zPvaakN2lM4VXvkZ07mr84NV+vFXD78kkRTxpSdbt+/KjHGrW+m4CCCXYJM+
OixFFheg1Igw5/Jv6ojMbjBq40OSksqEaz+anUaPrxqmPbgwSyQb7ONtAcBj56C76k66QFYQftKh
mAMOpdwDf6qHZxBkYW0e8+MpNZQdjsrhbpG/XuYeQqlesDXCI0hIMiU+3YFVXFioxZ73AWd3vPhL
AS6LCdi0H9K9OgRCgx1cVAuvVpnK5l7ejnYayQohiqZ+/VchMdw6neaN7adgBgpmSYMw/1FHAs2K
Zbg+m1c0ofNuWFasDhiAAWUxYMIbsH7VOxnGKPu+liXjpwqRUyHBKvjTARoPsyiDZdQOegrDDdnf
4NBhRoqAvE3NLzCgzdUGeDWVbSILQpztsLo7GrxgkxWiJXWiOs3ip60G22P23nNyOpoFf13b8Puj
1Vs1BzpELKZsw2s5BH8tm6rwA3dIfBjFrddpP0904fW5NKPWh0JD0VmGZx57dGa1ycTXL2lq/Q/2
eAkJ5Rk4N5/0lpkBp87jcY79QWZ720KOUm45nReJmTf1f8PnoPPut37uPXdIeUGX97F4hdDLbz+k
zmaUcCW/H4P31iTmGBeqdCuxtOaHclVA6bYISeB9xdQsleg4S9D2tIVN5dW+nY9v+KenPHvYkWYE
5H8W11G5A11dXVGF3AOFPzc4TnnElNK5BoZQ0n9Kfo0norEJKQv+4TS5e3ItqQuFa0u3qJ3J1BSP
seL/Lz0UbmiRcA5Sy5kx8kO6B5dmynHb6kUcZQkmS5yeC6Ke6WLdr7HbEZe8NxVM4O1Vc5N+jxNm
5a7t1OsOXaZhJ62Sht3Hwc1KydOTT4+0FxB5IPyVn1uU0rw49/K1N0Uc5Q/a4F5B+fHOsX2cid9t
/i/uZNqZ5BZzt4eLE37EJXy0U9PrEAvAqLeOzF04tH+ur8bUrTyi1qTFODDIMm9N1PNCWRLYY/41
f6b232/5axyU4vPY8eK5rBiS9DMB/pvukDO/wemzE76U71HYKwFr4WQI2HAxYj93AaQLYHuS92XJ
Z4sRy2SPbFflcbqLVhqS/wYI+LTTAVus4b+BL3aHZ57/qoA8++uzWahtSDYc9mkW/QBwyIpNy+uc
b5xrNfwRD1RMFA8+NkocgMrtDjiZ5elqoA9/2h380cKdlbF3mY3T6Uk7HOWH5TNalrw49yjF7mfg
u9RPOHkr6fSc395zApk526noSphlBXnGrwk5XaYpKRamqGG1dzpn6Uvj51xHZyxbpE0tVeoo9bpj
EhfThgryH3hFU8PHU0L8rNvgwFormURce/5vSct9eTdgj6izM42rrDsRTZR+GNNQTEoFTZrVhClK
vJzrp/+4eU9c/11Owgqje8jBtEpxDAr88w9Ewp7iKGy5S9/SyPHvXwB+gtu1QFDZZSHXJ2GyxnBx
/+CrqOedon1323/1ltHhOmOdLwEig2kBFDHl19dsIFFiXZZgM7jnARQIEIp5LQJnyMlIBmo9SVr6
xclo2wbFvmT+o07LQHRhRa6FJB7hI+SvzV/LY/klpOOUjK24LFrYfhBxWRJL5CLPpXWLMpPpnoRw
CYMP++cEw1qOVm5+74KQkPrXbEhwSJ5tVLuRNNzjrPmzk3us/U4QHOZ4NAmMFMNShWeo3nJdgY3u
mINNM9KKheoKvE3D9MYZF/KNnki84X6mPGeR4puomEDtDHpCxAoJcw6dYx8pps57b0jPDVXTxIJs
dgp8xz6rUkrZrP5FZH1Rw/QDwudzCcDh3RrqecOqW5l/uFrBBxgkMFCWysn6jdvO4AoJ60v/nG84
3Fngm8/fb7D7uSOaLZX+HW33UvnV+4uvI1hK6givxaLKftaXjlEoGjDqq5DlcJMQFfnwW6VoRWMj
kalL4Zq90W3a50e6lQ9vO1ORubkc7PLTQPS9gUT+YRZgHIRcM0cPr5+HFqWD78ZTA9InWbNc8q4z
DRcp97CII+wFskI5k/iK+S+zp5x+DId7iYMLdpJO6Ot/W0hnxHaTGNwmSYJVmLwOOBU5UYtDu9sK
Ko8URYt7uYYQiKlynyOo+qlbkOiazwl8b5diOjt3bOL9eNeb+g/lA9wdsLAmWSeIo3mGLqszybsJ
OdnA4Qr6NQtge/EQ3gnW9of7cHJKnGdRQl8IXybC7tnzeqO/anqwCmjXRxypd15WLjQR0VfmHLvr
UmugCvMPvt4Arf+Dxeo8FJIWGJODTbUsUDhQtXEnNlzZ/QWk1HH4GnwBeN9srQfHcDIL51tQUq4M
rGzpU/xVavW6cCl5LMUp26rAih5F/Z3kXysq+1CI72pmAZPaY92yBfN6wvja/qo3UUOnIdpCW0HM
KvtJCrOORaXM2bgaHkhQZ/eHHI9vZi7IK/PkHbBxxXl2q9ea1d/fiAlKF/+yxAoMM78XOTLpbvEL
H6BLP08sJsCLMhveEmac8CpTKOCYmHE4wyJRQdOwPr/V+Mc6Pw6SCgPDKRilBwzTKNABAfc3ScJ0
3LPfJAEPIZbQGa4WUjNNx9lwE8eHJoS0Kfj3lrxWXNPm8j5toO9Qtl39WRhWsgx16Z5kryzOLuS8
dS3J8nrWTF/3u0RFN4bfwGavrZXPEUn1yP7eU1JI9Rj8aKUQOrlGAwWfoU54klAS9GHfRcvwCGu6
Y04wRCCeMVxFgz+blaaiEmRRK+rMmMGL5btXkWDzQxgDwZDLdJcotV5OBNGj/o3jxY6Q9kmii1Km
RcPdbL699p06wg++GaBidtGY/riUhmOvg/783BcmBpKV24w+AhRcrYDcSpNgMnMEcGgiPoMH20Ot
F9TKLAZqTZT0vwhDb/rZ1UOarO7IMCBHZb8W9DceG6mZkVQMz113UH+BTKslaCwi1ogqKZAxuLgM
Saf8iGTHqZ4jaoDRVdW+b+gMX64tCfbHsPZtowgNGLhN2S0iYjKqtnJhiHj/mDM6XlMivACTTRAi
Nk2o/0/qHwn0s7YozEpglj3W790yxXeFWi2O77lA76qjvi+LsgSIQNQ1Nx/w0L56eQ0vGc1mEGXA
EBjVK4ByYKqE/G0PzIP1ReBGDBERTguix1y362e5PfWyuenXdZyyEfA8Wr3UNPR24L+PBoEh1Utb
YJy6lYUxQzaPVdBf04yQBFmowelkXxZBRfWJkiMtJSSYp6+XD8jWtZ/bchC+SwadNNiw+xnOiHa3
SElKfBRVlPawsZL0NiAGnkz8PQXVE8Hv1TETyXfayayBAnjT+ms+wEMg2hRrIMANHZRF6zguTaQ8
8CzMdek1ZTwHnWNDDKvZqqBVVr0D7KVMQGH4fCqGJ92p4m49FxRDwFSKdoAC8IPYi2x+VtAXF+9/
XQwhRb+Gj63q5Od3G+9KRY51A8SyiLt//3YhK2l6+/xm6NhAB2dybX96kcqkxgk1eQPomV0n/Lc1
TLb2aZEwIKLhD1xhVs4VQWWZVf1Jmm/z2CSs9uS3oMpgf5NiUrPnqqt96BVUPAfAn3hSpLQp7PRz
QH4Im6Zwgor8jFb+4PbcjzgSYekE3sMOhyeVRbICtxb5beYxDt7rLdr7TM8TBjH9wlQWJQPfl4/Y
cPEeoVOpGJjAbtyyrVyr15e29S6uMKj48W41JzRuEpZVVCODmGUxewQkrHK/MYC1f5oAl7NG75dD
LxnRbbhd5YNAXPZDMFkT19330youSTswROVimBaEhcCsRUdevdwXC7e9eyK+5VtSBq4Ujil6k3Uh
1yzMI2WRXnJNZwyVhC1IWm6YGTNLp9p1CFVBHX4tW/zfEBHFueDKCNpLwsxNidCgMPn/FDE62h1L
vbvAY2m2B6v8Rj8AcxEP30ZIBzDrsjtYmhGBvnmFFn7Gj2qCSjxepdp+kARWObsL+vloY8wcO+4e
cMGTZquv0keAsF9NMR0AsYj/cUEyGXlDNBLwZAGg49tZtfZyvMtwa0L3rMY7m2FeHaKyotLLacZp
xUEd/jnXNi+D2BLfHkoCcOIXoAnhwHai+K848KC63HCChLGfh0ornye3zLnnNHRLOXZPR3WVJwsq
KSkcu7GX+PTeqO0wUSB/etmK3Jesf3MXBkdI44tmnkdE8NVtMoqRvV/DzUAvGvv45zDGs54OMK1C
K/WUdSd9sg+xiBjqOO6M9nzFaxi2WK60isWCHJDglKMsvAqnaY4pN3cj/9naMVfdYOQ8aM3a099U
d4G63JrE19gvB1R9QGBVb/RD/50RsrlLNc+9TtApqSPvFd1tyPnBwEbbjLaWu0B6UqrKTOFAB6xZ
NFPZIbaMrkdVq3u+HZHKwKdilzJiYycCC7StpKbgqexMne+MULKEC3HxzKMhffCzPguhKm+3crKR
Pqz+WNWHWJGln3YVphMNk97pE+RyRaAvouSgS4rAstsrdSpe7AtPEE4vU0m2GO0UNiyrvayc6TCg
jOkhVnto9wCVyUsQBQ5WohuemnrOSAWQlKMENr1pAjj/kV2rPn1kPX1hdhIejy8HkMECoy3AQ74d
CiiFFRo5F1fSsbSgeUJ53WKxvExa/aKYCKkxP9tVWh3r48fJPzbE94X3eyDdI1ygXxuO/NwRSBf2
PsbT/S2LPJ3q4RWnWblac9s/3qlGxHyGjcw/dFMYnnE7Z3LibSW1DRVsxpzAaKRU+/qR462NFxPy
H54f6/z1gudOAps/cx7IAccdG54vYAlIiNLN+XQleTWEfTv0qEkt+RrDbr73BWqmw1JEBxhihKEC
lQ/lrytpy07LZ0AyZ6dDl63qGbOl+MKcQrdfbfd9dvKpO1YZEhRe8D2Su/ltNHpE8iQvx/Iplvpr
NcWsLMedMhP6BM4geSY+fyLsiKwI4XXUdOqLx1eRRFyJTmD1/kq34xJRXTyRVNumf2lThCSgZcEb
k9RmUu3EEFApYaW2OOO8b4seD1Qe8dJmz69rvSOBJ4fnIbM695q15YLU2LfcgwNROXMEu1X2GL6O
SDJDTIMnlyDH1UAkJzyDdy8ppn+c6OJe8mU/SfZdFtDSV+qhN0GbZP54pGQuA64p6aIwll3PLmPC
gDUb/f/BTd7y0xhsepo9MRJBiJPDhYIJic4K5WLmd78WayNv7fkDw00owWcR8iJWo4hp7oi1163w
uYUycVSo/LXJ06rHAJYTpC1AgKYz98FSqOkN48pogrIkh4tRE8T7iSoiMMhEbkS55CQapbGfN4JS
4emzv25Uppf/AKAf0cLITJw2O0Jm8qFYguHCLrr3WHkt/MgIqtxORlkamb79ZHD4u6dbeyxhAauF
sSpbcXohMl4xGlgOylfpnIQ0Hk/2NTfAwKPMz1LN0wsejztfLFMEm7HRGo1u3042ET9SsW/vOyeo
OuRP3DY2fbEVzADJAWtmpNRQAKPaA86LVVhARhT0FNHozXtDOsfzc9b9VwEkWkAAL2I3HXbb6bX+
PEbWcD7lrPPCHok55If5zVS5t2e72vXSzGUpRzJT2+xSd+Kzys6r7Y/Ma3qlB3WF0T/8yvcBh+d9
nDJHQLd6NfDM333SvIYj+MCSzGGf1cyMWeosNu30p8usZ7JGP7DPNFmW8lzMDGTIBSFSx+/2AbRh
kcA9vTE8OkPZqS79YutcZWPcLNUO7nrKdENny/DPUrX63zTEX1jyKeJ9ncyGUg7BsL3dwOOSdq4B
SuO8dmRTPxPpaMTZwPLwdhPrXl1Ectm0/Pc6pR3dQO7RC3g/vcmRyscUPbo5FoeLnUeR91hue9kp
WxZS636h3HMWuxSKdThFFI3FbZpUEMgwMjAkmuAUCzxChs8y33wAipllpRloWU+rujgOXHALN+f5
qeBKYBYdJoCRq1JYqNsDX4T3kskrSbzLfDeINTXeI00WmJ7sJFQ1d62jL2Iqp5oIPZ3gpjrQGOSl
n6lsbVc5PEJ5rOe5s8WQvWFCfYINrwXJPQVJk4B7/kEbyfBcHWxYjsuG4LyVAZI1qTGkmKE1umMr
Nbdc9F3RLIbXFcjbPsQdkqeqta9WhpeuMmGjUCkH+0d43Oq7fvF6kdb1o5YuP3jsC25Tz8/z5qLI
BsACPackF3e6pct2Q/w2iwyoyGlBb4hYs+PLdQIjprZO7kPuOC1BAWQtHFoYH2EzRe1jnMXY3Lj9
hHGbVACJF+exqdaQY4V8wPeJXxqlv3gzlt7W5uFzhwYwe90geR08SIv3r/+E5krjmOYR7WWBRDCK
Jt5C+49VUEPwK95P3Vt/1tPoaEy+GVSDUEna2QPLmuEry9w//BvO/PptQAO/MlIvSty5mm/LgDHG
VeOlYbKH0ul3/Se/cWoLcTHPEKuI4AnYQIxUCgQyvG3MQfpjD8XwdVSgdS6y6ULIAbzaIqRhq0Yb
pW6bHk5rjaedJhjB9BBkV/RksmUOK1T6l3Ffp/Uo9MKkuSNCRPrzwd7PNtNE4hkkAEHlvY1kYaOg
StavYYjxO3oxOPWKKmqQSr+UJvON7qylqWaqbm5mvoFGH4xxFDKpT+KhbP/wwvBUBM1ONf5S3bTr
wYuyIJvlpUEi3rEkuiFBuyL6Z3zH1w2eO7gFy6wZJgetGKWONbmWgQ6klmuK165AUGOlLdqLJxDy
OCVTX4QWrMv+xfycCxj+YkEDFT6K808BJcxBuX+OeiDdPdaah5yH5U+iKx8Hjiogbyl0o3/LMIR8
zvfPVa8NLd/gu4KdJRL65e8IFuPpFez9V7+CQwsrfjpuqX795ScBWU2A/jSfwCQc8ASI4TH+IQBF
Me99ljUwNGK3kG7iW5MEttolnOmmUZcdsyk6wJfKo3ymQx36N8g29wkCoJMGrHfanyj41MVmOg1o
9g7IuV7oC86V+X3QGgKV7dbBqSjbCzUSBEq0rsFqmZt0Si8GvbsfeX9uGinnvoZCVffg1VVvhbYt
396GXbPuDOJu/ZeEcHmYefsZcpaACMFP5HWBx3hM2EEu1rUjHqd0m/XUWuaL9n/SFG+HRAna3hUx
DvxbO7xEfy9rxIAZaEkfZhY2z8kHhi0XJI6+ZnaLEnAjxOns81PxiSbjtAnMJ88mXBsS4rC0cZzB
ZcbP6zFUnVgoTpa5TowtvveE8a+QtDzaPpNmo8w0By0z3RwX/JPKfDcD4odWUHtrF3qa0Kq4X2LE
T27wO/Jz3q0jhhcX6n5ut8CqWP37NfU0WunsyaQPZyApPk4ym+FwUvN3X1RTJ/SLQhDK8rV39UWB
bMoq3RcJMdaGXNvtLBIfq7NOCILiDI9tno4xMpa44aczGKXz9U69hfhVixRa7t/jmFins3p33ine
ykiFB1N6NhrqSBSzzPASV8M9tqoTfEr4Zz6LoxDVH3Y0EK8bv/3Km4ftcR2XtpOBxPfTuHoLSrTE
x3Pkqk2/Gg7wuoFWqkEtNGDrKM+rXMgZyS+tufUAmwfzEXviMGpKzDxwe+POtrO40jrJr5IjMpRK
YRhTycZHI82+ENUYmzNAT4V23ogk5l72MSoDtfW1MJcnrgIp5uw5Sr8XuFiiHnjx9MH9geaCTbjr
A5MhNDf7yrSPV3JnXsuxFPxoxNlwwRSigocjkdF3hSP/fuvInMSKYHD4LQXt94rH7X3fJ44j/TeG
2Qdf+8aHL5KOxPt9dRLqFGeSVId+AoVzVzhN7kOV+cJ629ld85egHV5i7SD/Uk6Osc3jbZx4B4JG
qypSwtiA661JIPQ7GuNp9uoloJ+eVYQ0OpI6AogfEhohkfhttc5HHlPkX/XSLoH9bMBq9KQnr3P6
6RO0Uy7XqL/ZgbAPIYZmqoXcbWqcRCfLDdjHDEvmb4qNSWuJZkYLhDvCA/CaQ0JYbhTTGFDXHID7
9UiEfiOMZBvQdMfK14Ubq8tp05FyJjdFUlO0NATXBZT79D9wIjOAzsUXdD5O5POi53Kqx8lkzWhA
7A1kT6We4J5kKXo+FAM1NRxoVJdDX3DH/iibNv6DplEGih/PQx4547QcTVBueVkQK8BPAtTYR819
gdp+sPGlEWx5/HobzWZ7KWoDTETveqVSHAqa6I7VaQCMnQs68M/klwNSmEqrcJfFNoHONcXDKNZU
dJkx47Wa8YObDzSZk64Ak0CuyHTf0fdzHYlxdu1Jboyof9LnKNGuTcv9N3PS/0t1Fg4/eTKoh+1V
HiIlhzQGk0hagu/2ytubKzohtsd1LN5jDZeFhXIbsxMiv3tbSwETck0UWzXLhorpHP/zf22IcghF
Gs6+pgAHKzI2jjmsr17zcSKmJsyWfSyKM4C2POZZdnyzbY4mcFGojlU6JfZRHzTI/zYUuRBFqeMb
ZPYGXy7tAJLd3O/hKQy92VycrTLULsI3Uoc1aZGfx7zyYt2AnVd0czWRbC2N7oSbA76epooyY8Lm
JMAoB+Zl/iZWgNFb0xA8XufoZTX6Xm+oLJyIOFKhvE1AAPG5TVMjUw92EVPhD2vAmxrCGnp+pPtA
z9DNwn2NM4k0a90nogSUbe1Lc7Kyn0vU+VTSoeB1NVo0d9HbfPVtyigJ7fGfoBgAGKHok6xpr7Yv
1HEz8JJL858oB6fBehLri9UX9p7yDzW39ph1PQX2gzNx6rr4pZwV+5LWj8V2anvU5W8a41gD9Kpd
owKLT74BpL3VaVnRkdQzGDMzfuk3BhecIy4g7Gs+faSe7Mf1V0h+Cp/UiezRUsCCTnyPWHiw+8Oa
eQ2EZLHsF9F9lpUO+0Ih4FqF17QJacN0h7lfDXJpC+zJEF6dOXF78aqCmegHImBzr1wh5K1rTcd+
RmZTTJ3fj0tr65fT9beVY913dSqXWdYUoFUwbW7079g0wC49Rf+E7lqs4SHS55kcdEQEVl8nAysX
McdkLgBEt1eqyNvZzkmoP03z1f9FA5P0m8Bc5srCnLnI2HzLJCxZa9dfLjcBfRKBCuSGNetWaxbi
grCavZ5I+6nHwPWDcGs0kIYr8/fiEFRqRpWL62DU1SLTXhyRwOQiXWakqk+GfuCOifwfg5K1EG/Z
z8N0mNOhOUHGov7T9w2c2P2TV713SgFK7TDpnr1WmFBz10+REgrKYVuQjdcc9uv1Rnni9farLNhx
To+cbjqC2VRkpBVVGRQ6fp9sKhZFnMXdh5EASXv5Nm+fx0tKADxs34x4/uDTMlhl5+NCmA5SrL6I
cereB4cYIZl3nP4DCIrgcZIO8gFZj+t+Nb0HOIc2xKDVlnEsvqO5zjE63zrAKsoEXvLbPLRHslsa
Qf0ulXZ91xezgjgvhwClgxZ54YjhOJXCvbD7HWPMYSJre9hvZt/hKZuoEefsUlbW3yzzs4a9kmNh
1RbK/gfdZHabocJD6fhbMPBMtR/HcYOedxnTSIYUftNMa6VEwqrM2UsMM+Krq5JJ7JOOhpSixxEq
0I7uNiR4ZkZiV4p0QGC0zJNS1R6ugTRgOyyl0ZcH/RWuPmxvDDXwuYNTAlL92QlBs2mdHS67RV8S
AOyhr38sb4uKAk7ite/j8uKEOVz1uDlmAJxPJdE+1N2RLcok2HtvfjBZbIRixQG6rorFJ93MuZpA
7ooRSRJC+5jmQG0i8dA4xJYnHD1JdnPBrgS8AgB73SvJXO8Fxq1ovka3ddlFZpOreNYoA5FkCk/e
g5tkETkTdZH77xkntEzUjK7AxnygVjzKbyXdi1rtPoXZIfAOLmgPgL8CdyFeElO8XunYHE26ZFWz
6EjR/LE524xQ3EPAcQOFA/KMmWjnm6/azGW+jxTH0ubzPWJdgYw9br4bxd19DDsek1YTQFFwL73+
Q4/f94VlcMUlRTovuwaAUK/bduXAcr+nyQ9j8oxhAR5h+Json7OH5sEyASWZxPaZ1XIN7KLpjcL1
X8bbyEI/0W8fsGbXRbeYnyDAFQGHZ9FuWVjEo0aV8awnUC6lovari5lI7xSNw4Zj/SRcg6GJQzzN
EPgqMoGpPfl+DytdtTl6cQ56878blLTAL4HxLKEI6CMxLy2LBxCWkw0UDD5ylxwheIn20gjIQkOB
rvOqjgHE6Kh2ACUgl9tueA2CRMR8CsWA2TIgfM/9rYZSBKVjICOTlvoH6co/LFvZxtCimoMMV1D/
5pw8iipxxsbBvaRzCVfVsbfyddlIu7+qB2tCehA426dOHrkxXaGJRngrhsNLn8H3m2d0V26g8jTf
NA+/naB8S09CagRh2fOV1+bJYrgaLGagcyaAXF5GV+Gn0VILs9uC8ipYUStXE//EM+e9JltMMZdS
b56k9zngWmPGGIM7nnzQptzNgPYHYRXHNDf6txi/wzlrpG6sO4VVcl98y6SbaX9z1xQcVNNb5ZFv
gQsuj353wzwc/isW66A7BHMzsKSIUaxVCU39P3E4Mn2kScvbCBX9VFW4d+hMXOuhmTEp/It7dhE6
k7ulkI1QiwojvDTRLAQXlaVyuUPgyGEyBTQSIkdN/n9hDcZG5roxc3dquB4MQaU6j0QGLGMiF3yP
jnRhu+iT2w9WKN9+7H/vJj7I2hsDEPgLYNR0UUlWdNIM3HwSx81zmD4nB5t8O9k5LSd9t9UeAU5H
gYZbJsfYuUP0J026B9dSV9Lp5RGGrczO9f/5jY7zyl6e/33lIxsoFW3RVQZC4OLs68Zv+yeNBqh8
s1Drq4nAHwG3kARYZKj4OvVUDZHU2eUN+irA1AMJNJWi2WGg6Rh/XF/POyQk63ZdrDN5zMNkR2g3
PLBPSxhzpuGYKpdUToQBc6aSof6jKjxE/syEK+WsEmU+wZ0C9m/faZw4mIZ89KVkz4HbWHCYaWCy
hQUVVj5DfkuQ3xjCOfQrYCi9QDUZiIimhhGH5/Dz+o7IX3SOZC2oSlqMM+Dhr4dC/5zRIfSGJAtE
Cmd6vzb3/IaZ1YMm0A+a4V8xmrIEw8YeeUz1z/R8SDkwNoyCintyW4S+kGiiCmjbeGvdFhM0e/bL
+YZFYAyww/w3/57D1c+YwhSocYXVnoDYotOybRtLXmnt31z/vQCdOGcb0UtEMLLjmFhhAtW4DYEs
Zd1P7CCaaZk52eX2Wg7KFysw1trnmTN4m4+GacQhNE7UGiyduCM++FDRuP6ew3rCgAycnx7negOF
2ugClHSZek5M82vWt9w1cHztqKy+SqrTy9IWgj+34JPZ+lpCan4m/a7+bwvOzIEpSMX1y0jCkE5h
3yFGwG7EhZ+UgmFVPA1ctyKPKsfZCgf/uuGWZH4QUWFxZNfULzNH6A/k5GYKwnLdmqKPfkEz8hme
geqanI7rLy8/Mx7jX/JrrBZBj7ybn/wSg1UaoYa9DzxNJ8Jy7ts4TodxcZV12xI6muKHz2zuf9vm
Q4X6UbvExZnE0WM3QvMOPq0Ni+9BEmkIcV4M1dYVIc1rCqxbhbBqXpKfTUmBrsv96UMHiEz59Siv
RXTRkxLam4T240kZQgOT1Ca6R8CBgxaYohUZ0Y96ZI8N749oFX+lLPOIMvhxYAO+W6a5luRbuHci
IVkIjNS4WLJ436SLZai4T9IDPhBX97nhJYupeC2pap5fny1Jcml7TvrwoqcCSMr6f9NJ02Z/TYpq
ZvEcxQChwRG6herTahsGCCH6O4+zf0hTgdRaiBUVaFjBdzSW3FbmP60S3SmvJuS9qgixSGWLtLYJ
6HSy5hMmlZzTnrPsAdjZS1yX1sj7RxZcYeNV9UaIP4tGtw16Fb4J9+v0TrdS8YrXE5lGYgJSNNjf
lnUBcAtthYrc05wdKvkk9tnlSYNdIzUDJx/6o40wWo7fiWZ0iZPQ0Y3LKnpuKY9Ti7FN+v2e3cq4
/Mit72OnG+VY9Iustsje5rnTOQvZ80cIBisnOSfEZYKvC9Wx2l5kbtAlLR1Q9iiS+sRKCsWg7j/T
WS9aobTeiHRNd6WySCRvgyqWNibgsrWrGYq5n01JwyBZQDIus42rv8480HTYq6CpYiJXgxjWGeo7
wNHsX7dOoJeoijmL1VKhz/I/qMpzgy9wf4aYuyTAcMA2CFKmNtC///F/BDx8tD/jRD9YDuS3a4jG
kidoF9unFAueA1yBShOewHHBRq3dKTX0LmsEVktnjlSqh/t1YP0M2az078pZXs/PHPSfzpQahu9+
ZQ4v4bTU4RwFRKtzBHX0nf32P2GR003VISdrR9xqblaYn7/Vz8NEw8lCVx2yH8oaFy1bCNS/UWh4
RR8BmyDNQ6nCdNSnWddoW9SRHYZX8fOzQ1JaSI4y8j31DUpzwE0GEx85dNYLXhN0CkkYWCqiYBss
heOcVjLo3dfJeehPgtbxdNxul2zk0ulKIlKKxajpO4zTPAyDm1wBig1kCKg+6LkCKXTc8ecSH6FA
b7ATlKkHBqyl5WAQNWil7+Fy6N2Gwl6YhsCMWszaSZWl8lxFjmrcoOgbgZbt3iFNjCLw3RgfOuHb
6xuqQXrUL2IASlDQlNCW4+7DCTH91Gm6lkcgHLn5W7l/agF/5ztgZ27cb66xgWaCWvgYqu0Ag2SW
QkH0TZRfddT/Leh7299VnCIR2MjpKJWCFvW1w3egAvdN+JWH+WQjruDN52dnznI5mWdBL5wQ8bS3
98qFzhrHTg4DR/vMZob1Crlc1xcrZlL/8lxMXTRoIqLt55dnTNEcTfUedbA8FzhtEO7PSNQsHK+s
CKW3phzUkiSi1vh5bVBJDZvUa0EKb52Ym/7lfiP2rHhWvrjwsj78HkNAde9ifBzUAct+Qsko6zdg
G3+4NSisrsL+6wULcFRvBNzJ9imckOQ2oEu3by8GXf0qs790ShKwjTaFy2dmtqcfCm0tEU9Vyi22
vusoNB1qdhY7FNyN5FxgJ+LbvfBNTgUEqOozYY0gHMy0LAIHx8Eywl9ingZ8MPkNUhTFqISMbAkn
jwJv6J3qF4goOv8USgj/H1aLzzHqaTidmpUilRgCKpBYPm40RgdNoOnD88oEhJZRysxZWaxppY31
e+FIOSvOYY0hLNXy9bA+yV/KMdroRl67bVx5VZcTdH1ODkbzQiq9vOOkfnUn5PidfSznkBp9QuW0
jWvyGtpVYDr3V/3kHw+umo7SWp/FBBG1XgNJdRhXuODfzpH/IOKmibxIywWuXyw0LkUMyUEMKed3
xYPY6uakslM3QRkqFxgTdhJwv+ZDltQhsyM92OuXXG/2hzBLs50kJoKKt9bBxcdgOZOVcxZic+Fk
pbhGz25ofajQuY0aI8PvERCsycQTGKZO3Y64kqa405FJzV/Kq9mpCyqostHucRwQESrdJqPbpQxq
/I1eQMzJSy6K2D0tjsye5KeYhMpoqjGpbIvPATrH6mSq6124g0grgTAYlxHRT6khkDlG/rqoQo8/
bUeVXx/JgMGZhIgw9eF6pedDe21osAFWCGn6wBFWvUAnUd9KfYguuMKzyJKQLuWZtbnlT5IPGLOp
AzFZXUGjTjKcMpeXDUmbEkv3nAJmrAk6JPRKwxbaPP9EEADBYXYLJR1P32pklx9iDVdLTitVUVsh
MixTS+kL1J7A/09R+JdthW77ykb3iTG1HT77ZNgjcmjeRbCsOsb4d7nX2U+Lz/rnyCDuxdhZgWaQ
N7OAoJ+kaqyZtNu5gkOhiRvFP48GTLiJe/hMVJk2DDjezUhoFUcjaE+VAMctt3NOOpoVvjwPWLeA
FbSPsRYe6gZr59vB7s/8+oZ+6Chy/GcmBV/4IPdr0kskzWSUKpYxE/6f6gRdiAshrnIUV8XsW+P+
WO96cpeauoUtW+G06wqlIBqRrv6E+uE3OT0My9HJ+/v1Dez22M5uJLBbdNF+QbN03GPIxWCmhdvI
rmlIkEAyO7xlNcFZGXKYgjF5hd2Fvf/CQ7HM5X42nLnFiNQsI6WWwvDVlOwrK10RHPFYnhDQmQRr
WENoMV6tPCmdLRJxKs6IN9lI0cr/nntaO0zNZ3LNa+jMufmRar0qKYEJ/7nFlmFUi3ZLG3FcHia1
lzMVA8Wnmkkh3CYJB/QxMraGTbPkilJijm+or/Sca+TH1RI9vUoWp7Dl1xBGzQGPJXtiW4nKYanw
p5KcI9mjdFA89k9R1ogWiXwlGbYCvlwuvCPGpTc/Tw7hBaf28pWouHhi2rMOGZb4/RQHO9JNGcO6
zCHeV/QoNjw6C/gzhU5FfHw5NWyNN4Nui+2p2Ycj6bnBtFi/4GHH1LIjhmUr0FOr7vMZP+dF5sKH
IU9Cvyk+z6ZptTWVK3c8C+PTlLTrFySQkwVnOpqRqknMsmj6tYX/KwSZNqaUo87+cn0gO2Oi3EsH
ihx6Hdx5QTKBrHf4efqDZeUgmk+Beaq7Lj3YqTCxlbw6CFfOsdtG+6wGBUC/eUFlNKmz64BFzZkL
Qnk8iyqgaPyJEGADt8y8enVRCmb34+JrnWZYp77QJRMhyZVHspAu9CFvDUqkexkweStXTKMfyrbx
ckiLbsQBCm/vP2eB4ejnfwkMC30D1yy8NbL5vR2i6X0GxkbEIQDlXMMceheFjxgvf8WB2uiSopaf
KynnD6s47zYBR4lNYKKuop5W8uyauiZNpQoECaoiXzNoAwVo+UmBqiS7n763gdZfWJUyA33to8AO
a40I8CWvDEMpXxwkhIXGa3CKYzJnJu9Zhe0pIeX19e6stxZkdk8HCNky++wjgQrdxTJbDjaT5QvV
68Ae5SJXESWe0k/u/D/yFmQOT0QK2qYpPYamNWAM2PDdXKHbPRod+ox5SVINncrpPBIjy9xoqQgq
uaVyTihYeLmXFiYTVpVPFSX9N9bctpoSlgjD7dBThX82wZknS22QHBoSCa3r9ZxNiniXDezEoRIU
1/B0aIeXaK1wegTU8Mq+NWRFNXqMzssW2wFo1KYAWNL0b51SJWjY3Sem97gPPQMUqpIAAvD3954J
F6GqZL0QcTMcXr9G4Z2CYAgc2XQPIwFrmrJvxNm48BWsycmls4oya1GOrwJSIMSG8jH6mTM9A+Yc
FyOI7/dJWMDyMPBD2twW26XzObnpGrdy53eSGK0Ul7moBwiYtd3Vmou+DSRoO9o5M6e+DccfyQYG
MUWMNOHui3EudIOR3/qNHOXCn9tZ4VzclZokgdFB/YeOU3jCWTs1mBq79VoDXKkg0NoZ53M9mFyb
ZAsBNoZATyDTy4lD/cBO0rkGvIln6daE6nW0pQAIxnJ+eppr/YcKuxqRQMV6DrA2mJ7oCuFoxVBD
19om5DotcfCyjl77EVnBveFew99ldyPKNw2T4z/N6KJMvIL/n89BM2BTHKmC3Fx/aItxYqfMULaB
F6VG2JwzPLCsBQmuBCotCv7GsGVhFYGBMYoeObgXMbTHyYz7Rl1zeqT+YZMm8IGBv1IvvGpbx18r
by8mF7BP+Laa8BoqM2iCQ/Jlmm6sTW2udQyYHmp8nEjUBtURhXgj9spKNrB8zezWQ1BhmGU9zM1j
sCPDOBwX7pMGH4kLKEvYasRhujgp2qJ5CA7I5YIzIqB6IebY1r75Bk43vaC15RvEeSWYUwgxpnRq
KqMqwh4/QGQuUXZ8rFrKwkYf9EYtijGQCyx7ZhoBoDlA6FNP/lPAt5fYzBFuRpvbWkSbX9AymfNY
6i6HUJsIvXjtySf6isTqk7twTohS0RhnM/Uaj6IU99kH4wb6q8ctVGv8LNLk0DWivHzuMi4Y5+Lo
a88SN1HTCtkcFYkPNt78FbTZAGK/Qq2IHcWVeYMUyiBQgkx6KR4TRvFyAMAsc/Dxauf1UhEFrwx8
TslowjvMKoghkCK0RaRyD1uP/wvQE5MJDV72TUG4vzro/7pGfYrYEeXviwJ4/KBqOcqbqW/pCwq9
jQejSj8Ymfc0w+gJmE+87rJdxqKl9HUtzKtZhnqTg75BOK4L+60Y4t1nHuzEit0zu4JaXcnJxZLW
x6y8mrd59J62yqiuq4Aw6HdLs27hM686lq64DjulWHCxsK0qFefNhyH5D9KT9U7WM1kn4PWgIrzw
zjT6h+i902WJ6w0KAfF1udcCNKT5258OMFPSkLtJegeZWTN8mND6WEgZ1sWDmqDrlX+MTGHkORDv
P+Q7RSnkjXRLY9xbZwN7NRnukpAiK/MnsU/ZWMJLgUgTePSACiWNbDXg7nU+Gb1qJ9sVkW9Jl46B
nr3XtCVispTWb4dH8OaaxXWwveVjD6GpzijutMTQYPjkydNGAzHxXonO7v6PuLSdatx3r99bhplh
0VuMKA08fXcr0Zr/UMUFQUYU2i7b6HAIAWYZyVQWy91hyeba1zwI701wbW17k54W5ejftMJqd7ud
W8aUNc8+hX4NOdQKGbJ3Rj8mRwe9L5Z2SuAAkU4AeRvUnCvD4GlfKuZLPsvxIs5SRhW/DCdmm+mh
agX9+o4YksS2zm2814x/U0E5aWHyYOwn7Vz0Z5VQCJ4dIFXl84McOm4QFx/nOcOhpFOqAk+GCW2O
QwzpUVB7fhYFWgoKjEDAftG8lPNvDXtGWjWG/S5R7FfeR9fy0UsT72oldpFJiggu8iOOA7mZVYxI
85ow1nTGBvBTT0kWfszSV2n3v6zF4RyOzEeJp4ToUBP/7Nf9/ys4/ifcjq4wEMPSGJf70AR+64nn
lTYHKKh91PQmOS8E8IZfKqpwiLCaELyY4NQqSrNuc7ImzBm8dt91UxY23dTSE4W1LHJciFmpklLl
uAKhtfTZ4xroUB3Bj+44xCnDH/AWm8xFY3vrl6yG2t6WQvMHdHdV/N0Qa5LSWkaKSIeF0yU9ZXGB
RAMxxGayTD+OYH5b3KnPCja1jAwpoH2HG72dZNQdMLKXqZ186Bwze5mibLWrDCF81V/mjz/x5Xf9
ITat9YesAgLhznzvWM9M+lywm9YgBSCfCUq3ursiTBXA8G0Q7/leaZM2XcMNN31QkAs8giPsy9mw
UANQ0marixlKO+aLx8/XhMBPF6eohM3p6+GI/izOdoqFtqKGzfoDLpbRP6+rBLSkeoYTgSjpeTz6
HlssUwAGzNl9Sk44BcLn6h5OQqHMfsdfVjX4+C9h+IzBCTQ6iCclL+NRFpxwTRpMoJYG1D9BV2Zg
x/OjtqmgvKFPEL7izqmkTvlSrvVjuAOhNFCIUMEeo6GUyTCuEJrD85exD2kNtLF0yOL6eGj9WW5p
wrRm6rSRcb29krVGdx8ZTFK+MfRXHsUmobzaeqe40fJevaN/y4ZWik1cKn9ZfPt2ND03n0xl0nk+
7Fvql3vpJFzzhp7W9/0pGJ6CR3dTZ5waNftbvXR8JAEoMO1n2w2Z6OfOJz2M5gzKwsP9+fXMWtPM
cdc69Pt+om3ZvKPAP1bx3d2c5t8VAcJYKeworV8wRQKNBMt1pqnfrAXS24dySisme+RVwy3hNGJ5
QcOep2kwIWzPvTgO6BqCWpWywFzzLnGrMhCEMQfubcvsyLO9oq0DblY/Nhu0/d6m3Gmq5fpKv3u4
TiHsuAwbCgzTh+aG1EO+FLItdaT0q3b4SukgEOoP2jIS7HSFffpGREB1Lfz/GoAFpPrZooMD/CJ/
3MhPKL5Amk0OG8PzFHfK6c7pnQWeh71Z6W7tX3vzSbyUMAulKWDB0Ia8aHFwwtSbOPVhUG7q9ALm
4ezVd0u7AHSvMVU87hHl0eAdqPJ97ZIiXUAD7Lc3WBMelRwRTcVaSGWF6i62ff75dkmp22ANsWVu
Heg20brZTU9PuLpbahZHfTuo54XYeIH5OqomppvvrXDOeQ1mnmnTKwiER3COzKcDfUiEXmiH20bp
iv+GtzOnSExZv2zbfUGdX7QK48uRGp4xmiuJRUTGkPLxsi6Jf0U7Noh1/5fDMe/Rhy200CbQ4q5M
MKWXvEb7W6+fkJlNGzZxUH5qTLPU5wJv9OUw7R+fOnNSjnxrT7EPdHV92nWjRRrSPdmJ5z7jV3i0
ggrNsFUFq279Kmgj1FohTtKK/mzpT7PN1vlh2DCYj4aupzfWzlG4OHx7ZI7S/UtYA0l4/7TmGxMi
D9fbz113KQJ9FglHFUpGKUOGujD7ccembn1mOKkxNHqlXowCdsb5+i8M9dHnqe1r/D6Ck8D3Y9bH
wVQnlhR0kOti95RJuL0h/hDsHvPAZ9jQ7WmxxhtsPhcmBDCcSQJwkOEUzpnmLtu30JtVNOjFgKNb
Ej8ciwKilbnsiYxZYJ7Ei+505oFAZu5WqDo9waad4cKOqCOuYw3dp/knBKqF0nms7P+e3bmeWFUu
KBepvhtgl3974uxke0cB/sKe01+g0/rQzXfKeiWuyeIJ5fKvpO0rHXx5VY0NNRN1x3dzK76ZFhvU
1EljHQlnS+F4SsTAJylpj0n/4whYn3kfmpuf3oMyQUeduFCkBpxlBReVMaPburdB9dlshX8PvFQI
eAHzw5zZ1h9+8MMy6Ka/iE5A5J8rTsZXn/N78wkeUqzKY4LLAV1wHnsoFP61YOUm56dnAS6AOCwo
dxY4nKjeeZxArmJpGgqRqa+DO1O8Ed/5wTq+BX8SuHKsAFm+seO6vc3ywmMSRp3nivFBlP6/3B+k
Elo2wPimOcOyTZ1D+XXLAr5omaKut+vcezjTnlYbCXZJlD40VR7cIGl9s5h8mc4LYUu9sOx1i/qS
qXFa3I3wYDbI96LnLIqk84woSUrG2+93cs3GSgxwM8sgR36r6FxGtztkO4xRPcj0dPal12ddQUCQ
sT9QjbPxqkLWDP/ll8ckHRsM64liOrESnzxcaz3Chdi7K7EV3byzsSGjIPZZoagWiokitLvTWfrH
JjYhebMBTtHxiRXjVXAauiCovEzy0LPFGmRYwqHGWRpbes5juYnzMDXejb2FxOPUI3PPq6M81G5I
g/H90LbRfUJMbwokiU/OTU5uqb1P6A7d60vaP2kb0JGoD5xl3Gn9r4pItoxic/exja5u2u7gvkXs
H1U/8xCFEN4+lm7LSIcxnYdr1SPPYvhPsPiSH+xvnCxGlipf+SWMD75rEcyt0RHXP1ZO+S+cbav+
M/pnViqKSQ/UtTC7vxu3K0n7jAp+r04YuM/12k3W++R8mBFApueDshdzxGOFE2lMHYMEbCsi3LPQ
VzBATIeIWzdbvxq6lGFu2SfF1yVoLnPKBbRrGhAxRAnTYhyz0SRycaIB0f22KWWyECzAK1ojCZX6
vWqLGAbdwJCcSvVNJbmrTvzeilG5HsyEzd401eFtdLM5UBfrqwgHyFyWOagvH5GeWeSUM8iu2j4G
Tg6dmRzmeuw4exIrgwWteiJYm13jRmGD/W1H8S7oU2h39uzwEyykKLQSVRFHeQw8Fm72yj125A3C
a8V+kmDRcQHegOXDz6irbJLAPjboFh82ql/HSJLQa/f6sRFDHHyo/9qPzPT2b2Tn7HRF4YDaXqlI
z7jsGPbQqMfWC7Nm+/AgfzyrpXyxLJdxA2XeOzZnxd3JR08GX/n1LhwBa//1XZKrBCdFqkgqV9Ea
ePVD8gwTNFNZz7oiqzSJgp+cyw7yvZg1idjZmxKP49GJU4I0syLhKMcxsdH3HL0Bh22UvkXCvT8a
iER5B3momYINSIyt0kiLWGd51xyJlfBVJTGGv4UtEpvYrKr8l2tNZFVJB5e8RxeFB41M9PRElBCu
5+lnZ6Fn02Yhoy72NGpceHRUI+cCMLZc+g47K2KYIP3nHDu25lFpE3LmQv0yVQ8yprXwMh8sXN3e
9ujxc7ZojcSZKNrsIJaYhvqP34fTbzdRldBybD+wryObqaEpNUNdmQk1wb/DqSW0L1X0e/0L7FlQ
NcAExRTXkUw9Ll6RPgvNdNv32ROu+xSSCkWMyK0ciiF1YJ7XreqYjFMVjOpvGUSrCjPWjjAqW0U5
pEyN1/EaplzIXEXZJ2sbDXK1KEhqIm3Gkyc/XdvsxERpvGwdd+uSQJScjDEWactArSgPvqXHlY/5
pkjvezUR2MaPkRsHS88woTW52Gl574bQ4nk2t91L1JenKmUU6tbL7BhOt0yjOtCDoNvevOBapD11
8JEmQLImlZoFP0Jv6HdKjbADZ/7yHgC+XFbDnQiun07xDK4+fxAx577N1OpwElRXEJ5ejaD16E4k
Gpfb/zR611UerT39vSxkx27s9GiE7/FemGQC6Yy3DmwM3OyaQnsjFjnTuV5Ec438To8uIJTyC9N8
GwxX6uWG58hhMUevT4TT3GqOfExIg26TFZrJXpGGp+c7dRrx305gvIxLJ1w6I0pxjFKybft/BfmL
+iphb6URBDPYaD0tlykQvGSqq76t5AJE4BCpAPM9pu/Uwmp7YC0BQ5l7V0rjbmGNK7fFkm9l100c
SUyATToZqX2I10dsibPBNm7MQqrMFpD6L99EDyW+H10g7+VLB6oTmbxk+DAP2CPcMHj9sOajpn/j
UYHwLszLOdbAuw9w2G9/h5tYB0tYFASg2ZaBcYAj6Ly0S42dxOrYWjSxiwoZpqq4VeocsuxYMrS2
6oJqwA+5+ZBXKuO7Tm2d4vEKExDqKa22Ujd/srUEwHvEJdBKpP0bqcfpl63jEVQqjp/USMMgENSo
ch0gaFAPYZs871sbux/NOdQ2feFINJgRhgSSYJFl6x2XQM6mHwAXDmdnoMVuNKaJxkrvuSmU1RdM
pHFexGjq3HLa2CJAraa8/+rmDnWJlKy2IgrYsIWTDFa3H9+LUpSDAKqsaLqMmgfj+rvxyVZbon8D
cPb6jJCuV/H2QAFMpWJcYw8JHOjtXTgrgDDiGCgaPH6U+xK30ovNld3U7BgDRTt+pj9VICqIDXdZ
OvWh8CdsBNg9zahhXZ/83F0Xm7zcVpzsHw/C82gQSTxaLfLrlcY7TkqLgCY13f3kB8xE1wVtUlJZ
HEsPaXvyC+we/hnWvgmJJ60/iPCQlssEdvpH7q5e4twmFHGpEL+th8vitOQGr8Y1JmnjZC6eanQS
R+BqPVQfzT1ZXiH1OeKZ1NePpXMUKq43mAIMSYo6kEV2Nvjabfau+il0vJUSwSmkkn1PZ+rMsuw5
UhuxFDp34PWAb25PgTv7tEt0/OAGOR7mM0B+XX3A4jmnAH1SrWeCujqRjA+yJDgQHZjtHsc6w6O9
KIcxb5BTNx16dcxqM9GXeyetQmZkQKLePrHuAPm7qrm+YduCwGpDR6h2pVkmKa6PudKNE+rRFQoj
l1M+TaDdKHgHt5qVT8ZbF9iwIph8s+CTVLbraMRCstitlsvbngfI3w5Fcewn89b0Q/SYgIxqnt5t
Xf7oJOGbLnNkWnG2e2VD3fmfeeOtSs08N5PaFbYClkirSoZNMzSiUnDJqinjAV44CZqbYbNJmEE2
sYJvBtHz9Arj5dPLgtV0wfzgbRB694XY/NMpLJkAvVmMdVVuyQX2Avjbps2sDWBAlb65+HSkzswG
/6u8tUvFSznYbnJeKc0wzTo3jKsIG4r9UV9uZQJJD9f/d8YGPwxH+bW64m5+8o9j0zemjztAgLO7
B0pGkLRSb3gzS16HufrDQQ+x3l7XfkkraBKAFKvhHTGeYmANDMqLKnGR/9LdJeQGQlrkjluXKv0p
i1OGZKHfR9gRBJ9C8vvBz+zNYSE/LfuS4ny8w9X8vfnmmPWHL8vm78HM/uvz/CHLER/HtkgTiq6e
o275i4t9/ozkStJEoSLq+u4f+X1UQdQDS6IJ3STOD6k23JjClehPqVkwmBZxKR7ocsXxLOiVkq+e
cEpVcC6Lgcd4ydeCXSCgE2iDD2xtntErVGY5T1Wf0ZrFzklSJ0bjcM9OWoRoFd/xpwi/fxDc6gys
834De4kqkAbVqGCtBv+LIQgmnNhq/Gl/f7ZU4fCBNLGJ5TvWH7G3Qe2ZxyavYHgCekE1lDSQwxzF
jfGnt8YEZR9mbFXZ64UWgWQ7ohFjaGvQu+AyWUCQZfx+2ROKUjhRBdoLw0/VenWNGZ2rS0b6PalP
QwgH6RxXezNIizNoXVR/WpnplJfCk0ek/BgPpiOiUtl3mPiME9W4sxAPrrx81hXlCOtncIkWQu3X
AMljMlD1mCjiAn9hJFvoG0uNG5uE7wSJE8NelT44uHMwqpBxDr/SqHLMv61C2WQqRmFJQpAlJAEv
S2FUJ7ZrDeYKMSYG/LkqkDczg13wnk1hwIpgd3gbtQGR72huWABGCo2fQrzFsrPV6EZ8Xegedd62
P00ebLdxrdunb6e3LGqTMaIAAFQErYSwTnM4NqaZ3rWXlBFhpcSZQDyoOp+MtrPWhNbob03jkV49
lGm+mLfqHtHqgzP+QmGY11GXIwHVl/J6oxvBH/9IfgC7jaPfn8/Hr+Y1BXQcGEFym/OuIdxuQr+5
tgsy8PiESMj7Z5zjSxigsAhT9+vJ3nJTbxzap5uTQ5VaYQKv+uu3vmUgMOfG6B3q5TfqRqiZR93U
/f6rqH4f1FY0gGwH7nhZDSwV4MQ4h+m4667tOnQltfF+0V9+Nudx/f64t4N4Yv1p7adTJHdeduvh
QgZRf3qax5i5SNyrClM4ypl7X4oVOxS/IYmeHtbYWh/kmtOSZSKRaLX2B3sqZ3Omih77Fc2eXGXx
sjzYHlN8frPAPcE5hgGfwllDhXdp3Uri3lSwYx6Ipz1iQcTFkf0f7pDB8H1EQlSJGC6Kpjkn74vm
C8vJZ/u3l1c57LTDahJ25u/fgLAOmtzO1WFbU+m3rclkRYSe2KvpAr5efo9DmCtg0b34i9YY4BGB
K8dtM/LWCE09EQb2S6SmP5UHAgX9d3mz6FCcoClQnSx15Stay8+Du7IpoeVZRURzIoV2+yXn1J9w
uI4z9F2ECaWvLPwjLnLpTD8vLN+PU2jBrMgx4en3ss9skxBDueeZ5WtGUxWeXIBtoel9QHHeikPl
9lRJUQYdN04cFq9ZVnpN2XORG4v7rH/Pc4Otf4V2jt6+8jlEjAnkWmTIW68KLaNlrCtgvMPdeoO1
/btHZrv7HsD3xTbKlho5qsvZZapLfrMfZcGUfrY26rohBKKsy8e8+7r3KGxMDgeMTP4fgCstmwMD
6X5CdKQCOc2GX2mFBUs57Wn1wc+G90h43ONJYkt8K3zepw0G+IUlRHVUt6eeepp7dz9zoElplbWX
q0xiDXbpcR00p+z/YSEqH11KIgxaeWCwIOCLguxStPWKIazEL1oeocqUXRjhtkWq5rs0NqnkO3RX
f1MFxLPJbpluXZnLruMaB6RM/fKxicjw4cYhMaZDMhloV2N0fTvG3TMIuB/YSEE7vpccpUnZJdbK
l5BG5erXX6bD/+PN89ICNkHFs0wOUWltQdV+el0+5ASYMP4S2L6HJDAtFGxA/18REJamD/9Poz0G
PTQeS7Sm+G0Lp7HncMhopXLddNp4LpLu9o1lArN8edQDV946vqooddhnOUdaaPl8OlDr1wDOkbTf
x1l9fLHLc6GLknKhum+zvhkIV7OgbOzIxTStDzL3mLlqf3/s2MCSZpRoRDpyzFUvJ0MW5XQ6bNy0
MY4ZLlcGHOI+rSkbTdPQZ0NtmaEJKZoJsxJHAdtg0lkf9d9tfmlsbPJNjLf7Slzh/BTR4eWoRW2k
q++So6sdFdT7OMsScCGtuaR3mNjZ2QGr39uT5LlqX+lot3Qg0mgBkX4ScTEX8ho8tvpqiYSeHl+w
6/wbn03e6jvKRp9aKGzuPlnf1PbeVHJAJ5t782HTuWVH1kgwUqpWXuDNSmhq6tvu96FxLEfQtyaS
dwnk1nxcny0oa375Ogk0Ga36euwBDEsT60K74/ewvEu3ToflFLLZL2um1PoQYdZ1mLtytF9s9VgO
HhFtXeDJGEcbYX8dHdGCUyIbQQry51TO2pxN+z3ooNppFzsOKlCJiSi9u9JifDVGjukSLnLj7cVH
qbXdUzng8HVXgFJlOysOwZ6SGa2HVwWh7ONS34ikzx2pku4we67X86HblNQtv9uh7iHEZprGt/y0
shlVbI8N1pfgvAnMGQABAkJxnlZkQangyUXU+oCrd/QfutM9cZYEzkLiVsPKwPM+R6L3w2l92pdO
dpkHbclYAOxhGFSWj1dc1PtHpCP/8ajPOZM5xDDksyETp9UfchsdoFaMjzNhvrfR430fh8GtTNE3
VzIWG3g+YUe8Owo95m6HQXDC6Q7+wnPX6dgN0t9RrUMblpEppTyYZ1zsYEwPEV5MGdHgoQhCrbBA
1aK/nlNFumtt9Wcuzv0CTVFZ+0PP7fq2rFoinskdVGiSuzTWjDvKww9bFVtH9SmbauIaHKacanfc
yJgSSI7wJZ5Xec6rbjLVa1i/ZX8nHG6J34QolXpRkNf6FQbYhk9obVFino+5sGbk6oHCGdEDDKMc
4A+4+6p7TM2DYrRtikoXs1INVuNe1AcWBKwa3/OkSqHkA/kgUtXuTdxSDZ1j/9iRaGKFE2Klj2h6
k6WKKl4uzXmnP2g4L0yhJgsNl9F5E7waY0GaRl91pGcava1oxMCWY04YPWG9CUXnFLm28MD4tGGe
i4dU931E9naPcLeKHm2jaUojnNjN5y7RYDTGlOlfd9cexIzCRVGw5SLbW89ofPVLU7aOYwwq0ss2
Bg/YwW7U+td4vFD5x9uhSekoU7OBEtX0PSIfDZI2oLaWCzUVCutKSnTm0PLUtsKrHdShg8PPdqh6
/QdVYwXT4LUy7gQOdC7+my1bxRBe1uq76y21YR5xtj8i54KTbFsindTHNmvpI59o0/YSeX6HNQid
/bUWN/xDWPlGxTKLO6MKKO2M3828dB8/B6/M3SHjj1LXc8b1Bl75Ibh64DFmC4tCV5VaMPlbZVBL
j1RzQSC91JUgi5u6Q1rAtZcl3D1RTodUp12CfZJpBvamSksK8bUH8K68z0lFXU4rGlwo51SOVSfA
YrsCqIJWuWlUWGXo7eOACn0EzVJbZzfbhxdmIq/FD2bdGwVmmoB74xPQhrNPUhEgKJywwjyCHiUf
LUp81lmBAE7jbNWS7Mno8QCQ8ukRQZ0iNoic759GU8orZGLa7AsRWE/KhsGSJYVFfEql+cMus6bM
UPgZ2honV53H5cNeGjbIaIO0mUI8fnQkEGm1I+qJhJ2IFLAxnpiVDv7WrMrgeyJqwC9yNGR9QG9u
4PrkcicBieYmWLHNd3tA48mLI+BwMBEnq27mG7uVDSdYDl6zIHBLvzsGWXMPzhQ46KmF/RrwaWTu
emzBDMWUn13f3k7PXsirzS5KKbfyi7dD5uDyuHKyCTVxj02gnR009c4t8INrGD/FIgdwyb1DEB5h
EWup76VxS+0CkEpv33ZBk07vOAzZ/EBO9V0GN9MlgY+JTL1/yWFYdRK7NJIDFULwU2rmtO8H/un8
O7F7XzjXlwo3QhNFiwX4FW35PvVANalHeWS96nNA/3W1nuXdQNx0j1tXHuvgSq/my4DnfS2bEqoy
pBPzEdKK08i/MghKn1BbAvY6Apc+sgQTlsL9o0aUW3RzIO1AGhP70sz6y00o8AwxKIvx19DsNKHK
P/5FqNo/XCnL80tSariwdRmFCGD+fsLAWLeuUNmIprykIEr5xgbB9WvroJ9Y9veWPByZvtpylHkv
ExLLH69VwhiZy8FFDGVLL8tt+d88tamiLIwrn16bDbe99bf1SxydmM+xSCMtDKJWZVabrMGpJcyv
XlYKzbGlYmqpa5nf7/OjNp8LOUdCP91hFc8qOK8hj+sSwuM5qJZ5B+/Ru1R1pZu/4J+s0KBtRzXO
/qiUvhSs2f5ds6TJ+XhWiarbSJnLy1LLb5zm9wgeaYjO54GFs5wWzCwJ2rQDcD9B61fJVF9fxSlT
9uaxVS0GHEJfCZIZbaIrnZB+HKi2ktXl0LUEXPezzJB3nNKDg/X7vIWciH28NQI/WQEFKBIFtqSi
zoQEyVNYVg6Z7h6h3mIMcQ1IvbvpQ/EtUxzFe5qYm8ZW4NibXKeacMDYqWOxPhhiSRiY306l+Ny6
9zX9DBWNtWFYc4Xil6R8hdxBwCcSnUMXr/+o9M3AKDkXBRYfJY+gX60GhKDtAeGLRPXN/xm3vzvu
jSedLwzIk+daK73Kr4ojJ1VYAdxVxhnZQi5iik7S6qEF5KPrfl8C0GLx8lwzhi8xhNrVm85xgwyp
g5EJ1K2glAKdJ/WvUB7+uUJfvY57MbFLapw6qpzxBYWgN370+oty7BjyAVxHozKtjrgasAUhq849
rGxRpYuWd9JRyZzFnQ2NVKx7GuFbg8dnxZ+J6bHWNfONC1qcfSOmdOWT2MezHVZ+JV2VVmC/Py8s
LyOaf/4L+Bq6MWQf4op094yhbi93TXp/cWEcB+wlOlAOOWbDinISnh+XmuX8B+GuzPIVeeNAf0IQ
fJv55cgZSSXEKMF0vozVuBu5xckgwdRWpZz2GwxQoEB/MKOyc6vwEfKDsswWSihpjfYqFpTtiuaU
KKYthqKrw6wcSwXN1wLXTSCSc0pcB/w884YdoD2C2ynt80epkKlpd7uojXLuUehjRvPEY3yaq4Q6
2qEA0pY411HdmSI7tE7wO8EvLYLpDDjddzlk7vL0ZS6eJk/WMssbHBvr/mBN+vttbN9bzT8V2wsS
b8pzqd0nA4HZnazYTxp8O7JlTHkORYjmKFyR7f2i2gkfonD08XhPBDdAE4YqMaSlpWWThpDuK86i
eT0XD7WZZZvY1/vu+kji+CoYIdiPDstTLbLqY/FyyAN8TqI5fqMIuIbecFpV0AVZ0fqxbV5uq/RQ
/hAr+ZyrVojIViecPfkmfWEO/+ktN0CymqAgWY6sibMy9G72OcGYAgRCx/tb54FhEepKGtYiJQZT
OK0Ttqq/1c+YEvHzysCqrglYkYoohNULuzd/ZmcVhw9fTmPvVuOlOT3Vuizgpm6dc2h9anujUVRI
HxOa2DA3ir8R9l/2HELtmhEmuaYfPjMjWduywFp/KBnUK5iEydfXaTqQSviIOK2PjNvHTq4MohTn
X38j8V/SPBpN/my/pSLTBhm/tjX4VbpuCNRciI1ZTI6cAwBQyRILc7mRjaEBWhkPzMRoj/DNtKzL
5tsDBXc8GUUpfORbEBrI6I5hPz+JZ97k/bTyv0luvHbupFwXCieSM3E049T7OHsr/LF0HgoAZpoe
lMcWjeIVZP825vjqSA1teOW95YHOIjQI/gHSqLUOO6T6ajijHoXFq6I3ni+7GB3gwDyLfS8OTb8A
KqCRxCSomjeSAb8SmK6lJSBmBLUlZ20yI2HBJgH+Bbbd4qm262LRLw7n0Cz0duA14stN7HWputoY
F1tcBz3/bEEYrna7hrluj9q8Zd55c9qNSVf9dqHY/tGrUqAhP2pYQVZQctDIHD0qp4i+joVf0tAK
K/dzKN4C1yhZGqnLTTreW7/IqI06eUo+GjHnuCefipMVLtV58NaVqz4CFDK7Y4o7Hf8+7SA3OZbM
3cTV+POmn1lpjIL1W5mPLIZu+kgf8tifNmOnKCGDFQBwYrTYTqUrQ63bfpebEF/mt+jVYMTvd4nR
lq8mIPdXDKEF4a/jdyqm9/62qBqwahdECDQ3lAKVA+HeVZnbqTPcHDogcFOnvebRUaBxNlU00f4w
qU1E5rOuGtsKfmO6P/d2znkX60A3RUj9D9nmTzlQunAQTbHgHdyHzPej8hEz8YEjY7lthj541hSO
l90Mx6TCo08Crr7p19g2wmuOWpPnQmGtmYDBh/1dwfuMwbFXdrLzi0JfbRr002BJzECc/Cg96Gl9
vvB7T06jpyLGdxKpL6I2ZvGcuBl8S23WRYAovJtszaKUvHHXWOiTYxt2LENwEgUpby9KPZetQ+JM
KRzHlwmUcGjXJoYwk07PuFEq4HqYOH0WM279Q+N3mXQdKcXFfoLhfQfkvzUc4kSwpeUqKnKt2Om4
4lP6UenNhefjJKWpYuR6bcpkc8NHfbVOW80RZoEg1Ot4p08eDhcdHqSLTEhwszY6JX/IyGrWuenj
zlR1JN0RrlnM0RmwZ/irIPM3TCCFwncXhfbUa9Q7bEn68VMXkejNIVWM9ehs8Pwl5YQJMf+LoHLh
oFrSNL8nOCOVXlAqcv8Bnrc3gWwXWYjT7CMufBbqEC4zOpdEyg9xhr/rA12Kpba8XgSymlArl9xJ
errfQsKIGzTQhKvw53Ov/yQQKtnOdXD/Zf/fdWpIUytGuKqzmsVNKNMK0ouIYi2h1tprPBKO6USR
kyHLe74i4MjEw1Gz8pBwWer3Wxxgax0hhNT01E9w2A0F6/wZyJFzExStj5ZzaM4uIq2aorLGY8UU
yU/MR36kZBNF2+aOhuAiVbaQxU478RdbCCzW2+cs9raxwI+N1AwA2XbSefX1Ptw67uTT9A4e1rDF
MQmHAeK/QswAjDaCu0VD5vgVvwEDr1x98qdwjcI5a1NQ9heJXglh0c3Tvf8wgTy+pVX5lR8O4eGV
2QtFwyeIAjeNvBpQq6Djt7mnHTRcXu9r/bvTs559UqZZs+Sm85VLAcwILongvDUFIm3oBXUCpZvx
h6KkTptKVyhjkMguslfy6skpKKPdbGNR0s0jLAgeeUDwZgl1XOwVHYQbTHszGIY2tonyHCUi2/ul
0V3GRhArqRwK+KlB+fspS2pzFLJVKcV20FiTGkQ3Y/KdvrMWpYuKEzPzk2CJ5f7fQQPvU2pXgPR5
gu1cqAjExSF8ba95JT3KamZIIGMZMvfSMOhjrJuyqozhfeEWak59LY4iUJJVsn+hQc6WwBl8qVUi
fNA5HpHIRrfskJV1/6BfrZwfwW7iX4T0K8wj13VsF6IuXexKpc/3XVlvRh7ATW082lkeeyYvAngt
DI3WfbS/deorI8h42TOhKPoHxZYwKuYVP8De0LJrxelr8Ml2IEYyeSqiE3pEe6arhMQl+TgLLeN+
q+lh0DBxqzwRcRfXLMABOYbtLFbTfyNW33OpFOpY03vxEjACyfS40cSOcjr1FTI5ULB0v2RorFNm
UyHT5XoJ6wd8DF41X290VYpM4koPNrX7gJkRCIP9+oK357sieSkMRjCKCf5Sl4qwe5Ipnba30X3x
BxsK3RXYguZ7+w9SiZjO5w96BIoqXCpoNdO7IHJk59MlzdKYzbe4s+yT76NrQiY9oGN4A3vt3hpX
MGwXhCxO2HLgKbhrOAY5yIF+pQS2ei68/neMcUj+IvcVtP6MjzVk8MUGlbYnLrVY3eFcQU2Gn3ir
O4IYHJCg6uulR13vInE57gKf93eYfvu9l5HbE98BpHUP0nOvoIcm6kkbHBjvKJeeNK74ZdWAyBa+
d+VO88vMlPrfq1e7SXqUkFqkfanTD7HafKqmFPncFi/yFMNJnskB1ceQYaCvSF5+DiMATzegJAfH
ZwBaKJaJzm/PThiSiCZPP4dsykYoy1ZrQ0OQnCIYcXMEyMVwrvKwjuglsb3TVcigbkiIRK4qgzTS
bJcy5DaD+sGirq3pt4/557MaGq+XD+spx4UPsb2cyG5r2zAfcXDZjoyGE70DGdJjoE2Ig78Sbcpt
USx0dE8hgFgNVIh92HGAl0BLsFLc9bdzFOWYzF2fVCo8QZRBRDCaCyYzSCFme+nP0l0GnY2sXp2j
kgKd8ouXeitkSYFjLu2qFglVW2KYNrNtK9fqNPQsrF/z6Y2gz2CnPamBuJ6TcGmCcyWKbqfNT02F
h5MECSNYGj5B5pLtoExn6p/P583TUGvA/mivpp6LeEfgB65InqXEveNqgtcc4AynW3xxN0rydnoN
zHN71Ldw+JAJi1r9AOMKWQEaJGonO/5OGkWAm+LZFzueCHdghhadCbKbhnlSKfU6/ZQ9wOFh+uB1
ga7RAYR8FGBaUUtk9saG1QTJ8K8ZyxpXMPk8UQL7ZyYoAUaHhsKhakzgpG3NWBqXZ95yKzCMHnzN
iflc3YlEGn+AiQMvBfTpScKapTLAydkBDgTRwfmRQUg1jBZkMf7HrVSbdbJs6VND1+UMHUpG8w+M
Fp/gFVu4wfrJ/2kqsPdKHtuy42FFi+jTwoRGdncgt367nQQYqruXvigSgxjU4jYxElSLKnqwRh//
z3jOXjthI5DJeYjBq0qcqb97R2iDFe+VE5R2QeuKMtRqr810JRr92bulRQ7KNN63C6ykLl+Jdugk
1rRrBcYE+QY/CnRvtHSkcZehPyjUl7WHvjy13NLFipTJGuRrP10HZ5GVJ1nWX2IJvVEUEk/reO40
hc0o/U5kn62SSmSIrMwwpwg+lBmK25/Vn8Gia8g22cZX7/qkqD9P7l6uFzRPOceDiWv3yuAzmE2I
fG9tuDx4osdhegfrAuS7vJkfKLvdweequmadNZrI5/tfV+tLCgrPcJf8bBJ8Uqx+QElSRT9n4H7r
3EVXFQrHVNmHqO53q9fQGAoh8uji8zaCM72p9Lgo9uyS5xC8aB6av16dzCztnJMc1qUYK84/3T+W
Thw8xKU/eX4NHgeosFlsQ3ajwFsVyVn7m7b89luxY6h4vJLj8wYUZzDIFfyfOXSN4TA6fu7o+1cM
8LuY0g6I2bMzKsEnFfYLheWnxPHDi/5/PQZxZHX+XpjBNxiUJEQzquDR5Qh6McwG59PP5ZBJgxui
vBSqRY5cmK5uNExIWKAGuGf3ukrw+d6ChH2Ss07sqEbqDSq5ALupVI1ZuBjKTQ0OuDO2nhnJWsE7
INWqjf+IkoRxhEStOqTrrR7GAXvRjvzMXVQbSBtW9eU+XW6q3x47bKndgP8GQEeceW9U7Hfq5GoF
X+XZcgGFY8P9GfZM1uUS/6dgiukTQGo7kx+GA/e/qQJvWBXbx0MKgCdfCdEH25s7dMwYA5yTctXC
+9ljOqg5DjYCm7SPxDveMJ7tRhVgxWRX//s8D5od7uOdYtO81EuAulKtxwO5vlSHzmi0A7Aa20n9
9VsnCK62QCmucOgRHHqg6JFys/YNZcTbFNmDRpHoXANJ5+MrzAfiT0SIabeOR+FzfL1ZmzDvhKer
xYg1Ze5AL9L4fC0dgSl21lAajy9hUf5p0pGwUlhPxQOF8A6EiRU6xt0w54pZizwFA29pgqtnVXOP
JGMs2WrHY9dxho6i4PIxAUzRPWcOztFCA0iJ/jBtwG/Kp8a6IJal/s3NL9CK1jgMpJHq8W9YzjlP
3sLXcHg2CKzHBQ3s2s1ufDFotbD9U6s6j8M1I4jMN5Xp3KIDkuS1daYdLYgCifYhaOaG8ULs9KSm
u0a/pV2AdOgvmCJWR7wEBrvBfLmTeYhIni4txX1X6tlVmMKieohdJ0nVnSKwOUgprwS/TqaLsDnx
sAD+sQ4M6/TIU88hI2etDhQYpuuRiAsGvlNmLiQfVEpyp1nn4N1KD9gxHPvMKsls0ZIrTznhjdS5
z3MTwOoMo+Gndg7VB6ciStCviYReT3wa8fJEt5h63GPSflXEVGxDiR/q8cBORmg9jgfFhUow9aue
oFl3v4vvzL+TnJO5oxJ1Jzg1c3hgicx8G+GO6lNNvDbKdJwW4WmDV0oGbos8Zgm4ZHX6Pv8nqJO+
jqzKf7ojxFI2LWLQeIW419mDeESvzW90Q19yEMNjcIHujxjFIXUcJEqNFQs4zVbD1GMPNoDR9liT
b0fFI6hNuoC7B3eIl/JRISr3sdmv89Dp1/tlljGixXtoh9UwW5uKIfR9gAl6VnSjBOl9epKybmWg
+KLtr8KuKPS8J1lCqylqAnD1AMlKu1u7L22C3nxSSIL6qyvZQP3eTT2yW6d7o8TYW8dMSEz2bT6B
7svoTO5ZflV+IKjwM1i6L8n6GnsYIwK6uFtuNI5abSAX1Ctr/uO7U92/JhGL0oHfSrw3D3W0YBby
QG5Yqg/6ASy+lfHnGslFUua6EUXDWG0+v1IX0pNMeIKRNRcO+fMxYqxJoQgvWl4YZhunZN0eRLQX
x8/OThs2tvxwITl96/xl0sIkQUtcNrlCRs5kdMsje1vMVorJnEOCZo3B6sBh1Wofm3avk0ABZs1E
hT3P2Sjuwu4R+JFQ9qQtr9F2MczbyRla92uORK48AH9GC6FCma6ES/YnoZRzqw2gaTPOfpiv/28i
344uVQAmYuciUPSvKx0DcPF2+Gso6VTeWyeN/jH3vVyXa4eoljHfgS6yW9PHLZ4ZhO6sPNXgWj3o
DzsXFfgyztXobpW3KSh5aWbJXSnqVP4RfP6Ik74bPPkuZMqKsvG3tko9uKJP5AjNUf3ajkv+QXTC
BxzxdtagccPtGQcIFdwQ1yjgGuUaZb/wXPGTJlzrH70YpiWSutrbascwXa0cerFIkOAYI+n/wxGK
dcRF4O7KYhuDd827HOCN+CrZ3M3szWW3otKDg9FewL4PpWhf2YuC7azK+EeK5d8BNoQ7+/kXXvrP
9MtAkWVQe6fPMAaUemVZRzLDUHhW1TMxoD2AS3YqCXjsAmcORDCYYcPJEC7SGw5B07GPuZYneVeP
vRwMuAmqXP3cJoe1gI/Y9KTdw/Z8XeHq035waub6R7b7L2PdoAp8v4nU0TBeKIPwsHn+4dZfGMPX
Ad/6r1mGCQRZHk1adIxOUK24gm9QUDIYvy9tEtlJ2AHVOIOI0CMbgljLMI5q3yPzk7LqGtOm5gzq
sXUtLu/IzPhmJWI777iASB77+RZoLjgNfSVDPEOp12324CdAnEzF+kx7WPgdrk2ZXZ4Ox1E13L8x
Sf8kQgBDlZbSHg7+SdA70q/thSsYT4pEBysg7b1VEynHIrBEDgdWkKTMTTPf2fytjdBCfEz/7lC8
fjgm4TrylUU3u+hzAjGSJVmvnplAG5xrfaWhzmAMnxwOG6K7x3DBj0VwiNzlfagQw7JKkms9LgmG
DQMFuiXyAn6PBSeM7ZtMfqkcIkn31ZEW7LmxaMnT41S8UDHImxFI117+yME6NkK93BL4MnOrCMNk
lf/UeyJnbLzKgx+UnT9hUk3nMIyCMHqUENNAmD4zr+tOwQo2Oy2pg/k6jwuzvk8F5zHridtTA7Cj
6SiXq5uuZRmWrmwNdQNmAtbJX8JUXRwpPtxCr+Sb0XY6evE55qBFR88WCz8TdXxzEK5alpodmmhI
1WwU0ogKp5kCNRmRfnES3NXS7OqWswrqNFI++EBCXD3bn5XyU4kB7u+vPkx8K+DIxqPfE3KgxARk
EbX1BcHi9Y7R2Z0S6wninUH4SNE3Hoo9kOYxHlfshRiZm1oc+g9z+UVauJKcHSOOU6LJktsTeYuL
ft0B3/Vr1NDmfEpZch/7F6TpQ1N10mYT4zwZrl6NE/A/oObPwd/qaAU+C1W0jT1hAl1jp4PkmrQG
vyJtlXKWdjxpG0ILC1Xk7D0Xr3/4N8IuguIhbb01WcTFW34Hp1lpc5/TW54DB6GSus7URpCXivHe
vOIKZBn2k+cZJREEP+fJYNXAz8rCLdxJ2AUjmbW2QdSCRHQOP14qP27/Zt38WWJeExog5kf6EJ4/
g11ka4up4A1hwtszeDvlKlqHsyd+6fO5BISyoAhc5/nlt8gpzFxYnq7ww5K/JlYYCfJ8jxxCfF5g
LatUVntrFBUsc8DIzVUDF7CFDp4qD5HdjwQP0cv/tjiHYZIDe3b02BiJtWPXXYeHPuMCt5fUTQCV
UIheg4qm4fOjXu3Vvsr+Mr3dBL3s4TJIZuhog5naNymD1GxC8fwQoDSPc94mjaZYUZSBET/CHClQ
n3Vbts/+tTck6dUU2o+infYZ+r5S63nCwy9EomUPlvSrUUoys5AoLWQrZ/sOuOobO28UQ9X02mc0
Xjac3Qqm9ABC9JZlISdXtyacUyOQRvCoJraayTWJjFt3A/2Ep9WoDl0enun2MPhzZ3kDEf9FQHQg
W2q1PN6Svf/e98K4DvmcJxBaGbmWQ0VxHiSHV5GaOvt52Veu6/eNjnY5Y4WCwJ10YiyYGFM0e49+
4ucns5o/I+jB/fQz7h1PKFsmsoIv2oPlTnvcGVUkXLHmt6/8dem4VWrCqrsc4bElB1ToiTjR9+sv
2AvRKeFpmNuyFDMjrDMyXLWDccX0F06iguXRUPSdT+alHoUsUGy/q8j8WhcVCVHcT+fdVcMy1GJB
3e3Y7UzC3Hm/kCm1XUk5MVF7x9gXmqO2Ze/+AMYu0QulwPEMo9/qSEpgIKJwvIchFdQgLmc6JoRT
9o7AXX/Ma5ARE/gyJXYFv0NDMiYNJ+ZTcEYg+VhBIbLVJaXDXTbZe0wzKDIIC01R0HksYoOi9Www
Zp+mRtdL4wVAfr/u2W+gjvUJCGZhLcDABXC5oqjQfuGT8jAxYeJjS2Hzt/MIdxSfzA1E+Zxpz43d
aucctD9KuPBH1lr6lXkPbqHsD5uGMG8RCcNJB0OOx+l+LW4hT2DSsXI16pOM5N9lT8OPmvPyTixY
5ghe46KEfOHnuttceNIQG1+SM1eWyd6ufjl7NIWbLJxtke1R+5IWXd19vRayLtobocWCyYKsATpQ
/CPtkY5+TtOIqErq4sGg0aMfZ2sJwfZQiQeqKNv0QnIDggeYMARrvHSaiV6YymCFfn3dNC795te/
k60QbSP7rjBKtBiLVgbZdfStyTlETgF6TLKgXzd3RHtpc2XPfbkmij/Vh2/wA0EaQ6ubUqi75ds/
Tdcqr91WcweFGzalPF1uTJkqRtndNbnh83ngSXq7WvJI/a0n7HP9TLYk9xjb79ym/f2Qy1vq/0cr
qOnjIKhafATm3jZMVDBaGj51kLlLhaQIOXR5bo5HZAJibVELl/6fZUhyTyKgxl0zT53yTgEWAwOr
Us2QaY+e2sY6iyM1VDrDos6mhO++9odfkSZ4YVGnV+/KLfHetDBKa09rIljhv+9Vcj13uFrWXZL1
9gcuue3ssvBTTmG0Ttjq5bt2rIEKS+M1TaSrwv3Z9D0wlijJLhd3deCs/DYtFmFGrU1YhV6LUySb
EpfNFzUxDOgnn8mCXpraYJ9Sjd8YHo4fSy/6HYwg7h+lsFhFtwplcwGnvytEIpgr8cpeMdFSLvZH
eBaFjlZaNSBw+8Up+STu5+4Ym/gAE8jmXUnJmm9lEas67Ei5Sx3xJT0l5xgF2pMwfOaTSg/I2qPZ
W/amjV+ine57yf+ymWdW29QgWIeD4n1HT86kjxZZeMPrACQAW8Cmh0rOLCiIei90YLMSUI3Q85Hr
F/pvM5EdDXRjf7zeT4rvsSv8HIF1HsbHhzWifcl9GHN/SkrP2QtuXpa30nXoKGJ9LNBUdj2+gUVi
aQtwS9MapYFs/0Wb7LqWX2SlMBUwulRwD0dMk8e8tWbSi2KRjQyKq/6ys99AzfAJ2iZMweXeqLtG
E7sVL5xpw7HtDrjSSMJnDYctufjssj+fuqpGJp6yepvklgZYyudXXgZE9ALD+E7MdrxjGOM11Nx0
oYrqIr5pvq68HxfTZHIRmMO2dvjXmgV7ybARdTUo1WCoKAsiZgEH6v7z6FyrQmKZyCZz7lfMPwa3
tCEygQpXiG7oYrHtjivBOx80vpXyfi4xheBecwSZG6/LDmjixlzyGcQYOrtdk5p5OW8VRnGvwUSB
yKozMkXMIFedFv951sjGegDwyfKkpASK07I5ga3VmYaFRJxb7IIAS+xBY2htWsQSyWCOlwUpJW22
/a0zY99nUgXC6TX+veWG04W8H/7sFopq6hiEuMEZzx0o1hkmlYr6tnBqi5eU8ZHWtve9X0maAExB
FP4Y1yYhsogbB+nWdNZO9RFZfuas7pjqXsW/BNHSI9tyetQBSnzv3USy5ZkNWCVkez31s+qyUvhA
ugqrxdNZAuGu3gYdwILZlm2wNtMmS2XQwtfgB2vMGqfE1KKYbLPZFAVuWRuH0sT5RmQUz2cX0bQa
IxY94+l3HI4ObHfO/f2pz39CPWaA3X/mO0sO7akxQx0K0PCw3heHvkE0YjITSlMRIZkMuHqSRY7v
PmEXv1rJ0c4g1mYWFONLEXaf835VmCt0lJjaWj5e4u0uD+PVievQ8SyjOjF93g7Ae6/z4VJQZGeb
hxKX7RIcDL5xzPwDI6/dtCCbcUqp+et0IkkAM85wAgPSgyBExWzj56koQfyyzgCtmYYSoFOMXMWO
t9ScyeL8B4uBoqU8hYa2K1szUua5SSOfLnBHWjyX+btNBFsFB5M02ATjWkAuJJ4Uopr4ivEn0A/T
2JVIcI/QnK5Nd5IchObkoPkmUPyKP1ZcSDeW0cuIv4vdL5S+SwgsxA55TF8AWV1QoI2X077bAsKA
RtcCdgJzW4xxEvnpxsEJ2TO/AHC1vKytK/aG+Mt8hWw4J5fQzIAL77kBFXUCdQBiw3aYvP/bBg2Z
y71x2051L2wS8x7SeDyz9X1lbtnBgvfBeAmOob7cdYW9jiirhgY8ABB6AaxF5DxwjqxDMMa4L/AP
+coAoShiPyXPS7LebVbA7VmwOsSqWTBXcR65kX5eSjZ1keFPdV9TuDmFnh6MMzBlsP6r7Bjiwn6q
UoNzFNpsp0gWFdwPc3CnIk4IBEBaFKCmpUTsnaucbRkT9wWKDIA6G0wAvTGN4oqAsbRsdlJ3DMFC
8KHcX3IulUkOePvkAzxe2q0BiiYu7LsuHskdRq/E18oLDhe65JvOq/5G9Y0CWjBEUge2YVDB/mzY
aCcN2BDTPEwQuotEQgNsKgoeIjMQ0Wb70xMtFvFDww3Z30vKTKF3rLWyvXP6HUozev9t3RVjpwpM
LbL1eQlaEaBkM3HkSQqJk49ZEwjx52Fhozyv2n65LJlNDiO8HJMYdfZSOQNHmFec1q8xdy/9wccK
nIyJ38WyqwOdqiEHiZ2OzsSOomEYLOYwIbX1M3JRQAtc6rPRxfjN6Qq4glESIdmIKaLvjeshHOyP
d9O2hd7LJjuRkjXDnO/mvsZ2qqPuR+t6z3qsofy4iz/KlYhE4/zsitUZ2NJItq/dzqb+AiW8BExR
3lXb8m5qgqMU1DkBwIkVSXGExZ2UQLz5a24UyD+iE4+k0qdzPJqjfOTAjXJG0FQ8eUomjVF0z8Wl
3I9chXHLAULBvdfdF5ascLpcs3Hkwt0jfHVLl0is0pI19+0AQiHwkrl15JVRHwHbGAiOBRDs2ktb
uV+SthVMUabTZ3e3dPlgAGmljm5hCBT5ozqslXzxSuyy4sA34Y/F75seyEmKlXG6CzAoTMo8DWK7
646gQsShPI/5lGALsYN5ekpJ1j4FeHFpGeVNuTnJBC2widYZJ+OZi5RCncC3rQufEskKwoeZq6GL
neECzu0skEygBJm6HrbBk8otyJsD9DKmhgCzdwqdsGhct7NEKVojNXd1F16bWxMP80Vwd/ZKduco
vlo/a5afseH2HHIZUE0u7Wt+oQRPx6fAbr4z1mYStki6jCQljWmSjhq522nzYFNcfNx60o7yn9+y
ZQiKxQhAKpmhJw5MmrA5Ijd89aafBWf+ohN4eIRDaiQd6aBgt6e1xv7MaSt0gCorskA8EA98fvEq
VrqF/qZfjqtpUCiIt0tw7WsHgJAVrHDpyrhHKUTE91Wk3FEnjq0BXccwU1o6DgABqiJ3pi6TSywB
x+037rk1ezE8gFJapOVV220Z6J0T7m+1qNQ7kw2mZBXIOs8NOokLSHA7JiKrLqFOdmooUNGxNgyQ
ODCMYYAPq2NxV5xltpbMe1sg2vXxIvjtOcIwV31qbeGIbMAN5NPffh+wpAUDSDcjvWr/HUASoxzH
EeTHX3x4qnKbXiWBOD1gnSEjhcHIF+eL+omnPJbEn3+OcZM8TsMbdTeVHZQeBVjw9d40DcI0rM97
JUpr9400hW+3TPCbdpP4z59g6ht0wuR2Ex5B5SvmxGyg5jmky7Uy7eLmn5+ZM2mZTWVbzB+4TDkE
3w3nGiacPrrBDxswE7tlZTt+pRZGHAKDK2Oy7e6XXYqYuGQcW5/jDx+2XiiKLOgdNUvqOIJWPGSf
QXKOr7CzDSSuUfJrEKcatXCcWg7CQdV/CHl8CXrhwM6VTCqYf76LQh+4dhJaN/xvdEIfVlSgSYPU
NSDdw9SySqWQcXhVIFyjwMmEiPD3VFFXT2UPOtxnyNihjeeiERg0AHliGpJ7KOGYZTaq1j3x+AlX
UxYXl8EVyUJbdMje4NsY88tmtitXz0UWfuF8Qlqjt2SoePHomx+L+9EILnHBdPgzT40GZC7GgeMK
LPriZwoE4fEKxbFesIvxCaVmEQLrKhZvOvj9KcAcyy1FdolEDYYdj2ybhJG3sO7nfsTXinhWDPwp
EcoKufg5XTEBdrDloGawgVkH+B93lfKTZ3Pgy/afb/BL/MnQ4ZjdUMSHlUSxRMGPiyxtV3N+R0dr
ppPPSWbtIPe8gormzwSVUlPspqgh9fa/lXm7Svd3UVzib+x/mt+JrqZZ1GjQcFe9X31gC2WfGjwk
L14if+2hd0EikdR0BEembEq0nrdlMl1sTioHNO/co8hMnnx/2CEHNGoeKF+/0mU+mWoY8lemVWo9
sZT0JdYw9IdYAhH45cdRHyfyrVYziMjQdTvd7PCQjDdZTKt2cvKuqrBzDNpfi1MUH6v7F/5gRAcm
S7InTvbD0s23wtIS0aVh9pMryKwPwG3fw0Xvz0VFLtlZPOZfdUsd92SOYDXdh33G99Hq7czSSs29
ewE2q2i7hxspMmXtnrYqaJuNHY0w/bqI/RfWZquG77x38wAfLXMl4NhY211VCunLlH2uVX3cWjSc
d682yDBUWAcHRCgMAbQB7I6UoWjRgDvlE4JOZzvoVAMy2r1izaLEto+NUvJBV1DjcafNRi7hn4Aw
/8HXyr8aAF/le8CenoKGcF9UR4kMArsB5TEaKk6fF3JwVidvPnhD7Ywmcn94zXpLSp9ZJJs1YeTE
3Hsg32hDiTx5X2PmmKA6O93FJYD+i+bjAhdVG0MEct04K9/ioC4SNgj4GU7vynijb7/CPp9lkXHb
pTblOvTsFWXs+VwS40BQmdzFcFCfT2Ix4Wx3p/16QeUajivhZ2aedTFbXjep4OzvTCd+bNXwoMIX
lQ+8raFKYmRjY8BGZ0bSxzo1V1zFzg/3ivhqbbLM1nvZHFxS2ghDyLEdEgraDRHBiXqy/vBZAivt
kIxqsXJg1nhCIgT7Eqb9Q+lwKg+xJqZu95yCW9XlyKIEF1r6wzSXay45meiJRVVbgk6F2e+0Mwk7
8KgSM2IhVQSvpruGdOXbVRo2F+VslH+6VgceEb3t38ibjt2I0YLmDIP2xoNjmCu7rpPUMhdeoAzM
wMm9n5hpbcZSsFH/urqu+fxBw8ZSYyIT40te0agvr044oznBzowHWIx17UAhRWoupMr6mzMzi4Qk
an8BtZlOXxuoXb/Rd2qW53sBXnQMsSIfkFML2yo34kUgJ84Sm1DrvSZEtw2+cV/Oh7I5FKhOgSNB
ADTUQz9wnTMYjKVk+eWOAFMdhxXv4BIzC+OVIYxLpPTuFHlcZzMiESIwZSSnucJ6/B0HvjQd17/c
P9FwZF8aYIdINE4UY0OJG/wzIwS2t2GsXKz7Fe2EBW4Rng4qsgpIh1NBTf3zTAfjaPh1zVmjPw2a
n1/1DlfpQYPoj63jh/uYv22lTRgwoMWaEQjKY0kER9WopwJqtcsxSMA526+ZNkLi2eeELnjSrQyO
lJ4RWvwUk3Ex/e38aNhYVa86LQlMx4uNcjbSM47o1yNiMLPKFYAnKcNs0uMTRScokTovxTl3x1q6
VE7p7qNAsZj3vU42xdA3ag+UrFZ2vFCoA0Ua0uQivNmXxIJVEoQqDVfqPCUSt4TgfeXkyRJ36ipv
+QumGfUcEl/qTMnY6QUG/Cc473hvjYrohIOX3gGgyZCbSKrEG0UXF3XctNnIdIj4D2Np1whgWTLB
UTG+t62aAgRI2WwXHH1IGPEkq4+hAkfQRENakNcUlpLhhgp5r3sYCn7YRnrrfkX3Qcf+FXiSVsbw
R+8nTQaFjdwSGieulysZcfC/42NqQ5CzYirCLooaviAdj7WrQh0U33fuSnOA8R4OtH3fLJwmemko
Juarrfro/ExfNOSeZdocL5fjbi23zqonPIpK5SSA3DzGDXg+/49g3L6IvMFekK6Mfs4SjqGUHVop
yEKyhCm+6HS97uOoNdrk+39sikh7k2hk2wwFHFO1VXsseoJItY7a2SLY1Yjzzf9GMm5QGaf2ZyLs
IKQdMPabmo/benvbcut1sbNcdSj166fkLlolaH6yEawH4q+whHLo3+LfT7JOVjDEKR2fSwCLf2I2
CHI/cWoquEpBc4Tg/ShqFTkTd3sdAeJQNyIGAnpgwp6iICGIJ7svURlnXoyuiNLQWQY1RH450wCZ
WGdTXtNIPJs0+/qh2NjDxX9U8XvQzsSgOzlCbmS7ybi0gWgVpF+koDIdaFoZzNq5Qs34W3e/5+K5
gVWc7g5t9NA4vcPXwh8NVJEUPsf6BHOmnav7eG0WsXp/yeSUOJS/8z2LGwbQq4tgrsKJUrr4QkVF
Eavz2gB0FZz9GyrQTBi1i1w+jm887gIfXl9vAvtpamUtriBgaSsoE63PySLtLeIRZHYzAKOvLzO+
/D/uI3Lu4LA+CvYuvnnIF0er4CWoopBU4hlpcYjsELMQI34e7hCVuFnfEPsOSO3IXUDrN0/KmD1S
CDiAKifoxGVAb7HpWnoOqng9Tgj+NTxo4Cwg/sEdrFKFXWCogeQUh3QyGDq7l2y9iSlWHmhm747w
RXCCtaXivCI9AyTdT2eEC70s/MyzIvWZI1m1mUaHsfNECKkCfaPFS/lopODK/7ZYWIMRUEkEpn1Q
fSuvseVN9bZJcVP2suo6upriIFZEtxs0Bi3L34BW/bLyVBo8NNnNDD8XaGkrqqZ4yas2v3VMrf/y
n1dDzDfRMuVBtk4PizoMVPYjkYnd+PsqS9qI+c1VB5tl14G4ibmaCXdPExIHF5W9/AYDWdgfJGGE
hDvV54wIm9RUJwdlkxWCMzF4C+0pt/zf122GGrbk3aU/HZmICRE90RPvw1+s1S6FHd+7vUlU9LIG
iuT73LNQz9PlgLZwUR8L9BHtt1t3FrDOtcQyR2dqbdyKXeML2UWOXl78aM2dI4N/iKAR7R1RmdTW
2y4/tcX0N3u9uiILCrQtqZGREYHNioFX9Wr3lBXj0TclWVYZJ/3iFjaqOkMvRWdb7q0O1aAOPg0K
5h1LQ9bqjpp22f5cNjYVevoP7S17yHA5VXYmTPn/Gn3rSycakn1KAisjVqF/j48MKW60eF7c/k1o
R20PhbrJVgCQPUq5vl8jjUb5hYaqVLzOzRTgYiccrUAHb7Ol1ek6IfxBlHyVQiUn+5U6UYK6/yPS
JpPgs38mcXEcWIhVc1z1UHDLKuoIG36jUGRl0JiokiDU2oGtrXIq05nkGjY4a7U6TOl5LzdaQ/Ek
0EQSbXy3zhGiHmNzggXmcO0A1zfTPYFVgWmhxLOXsjC3aAUV9lGYcYR+4zbziHg+2dqmc08jgK/z
aeji6UumAvXKhwpUxdMpIYPoorRPmv9BpnAnjLm9YjuqHzP/NtPvEXPWnV+qGLL/icEPv0vs1Tal
CvER35KfHrpakj9dfaGAX5GbJUOS8iFmS3FWNjYbc2733CffhTFx6AjZzQDnlsShCC1zHtPaLeg2
El9b5lkdFDSHqV0f8koMaICW0UnmNjrfijfEZ8UrM5AcDevu0qPxcpsE8IkdSYZdppcjZ828Y7Ah
QHpZNNM+uxZ0p1+rY0wiTYdIGq2/ibkXPa1tgyzVynBEJHpx3bx+rHPbPgOy0L3hLKNFPnyw7Qmn
DkWvuLqlko3/L2jHKHHTKm6Y4mrWrJOgga3Pw4zjd1/a4dsu1wu2Dxry7IwrY2kM+9WxyPIFL+ND
v4Md1Ja+7U0FoxN2022pjrCfbzgFyzLRRJBsyFDtwH0UJlOX76uIwtWPoYdDiaLMVv51vCsclj20
WFkAkmqNq7VQu/LkEFHI57qrCmm6HBeDVxFpGR8O4e2iX57OjjPEmvp2TEeu8xevmECnWo+V6fDH
XbYTOF5re3vnX7MdggwEvnRmrpKJs99MDQl7WPbyClB+ubzE+XIeMh2ZUt+SOpgHKLRsB7tSO4op
VWwpHOPtSnuE2CXqeiRXxN3KldBx8bdIuXXCZUqOKfTfGRg/AW81YZOe05cfaGfRSPjHiJvmdHL8
ny8PT6/x+A3gQv5TQ0YYd2Uuiv4lB7iEUMBI8i87zkmza4jqh6Tya+zhKVsguYDtn14zLZMdxUOH
RPPlYjtI+ckGeH78EraGyjL349BQk1ENxGLDRFavRwENvV7FmAe/xuzgfEAZjqsLnxARJnRPn0gv
SNShSITSHjaW0RA0chWXO22YX2pRHuzMJFkHf+EeL1rLqrKCftKIc7zeRuzm0Nvy278gX1lEFZH4
ljxadXoZJCIWBsu2NAn62Q3868SSNxcqQtMyyahKXH/O6wyLvrjt9PbitsC4HBxp+FFDrREoo1j8
4rzsG1Y/u7zuPOMjRi2mkSMjyfwUAPJbeZmmYHKRiQ2GvlPNzKW0fp/4yNvgu3uXeXIj2tWQihbg
RPvkIdTQLE3aOFEoAyG2jtfmNYM5XeDqtH+xyd5c2ZFxMermn63EgRK7r1rMpXC9zf/XZwucGVKo
bV/0NtOT2pC6OlzftJO0OCNxPMCBiwp7N7rwDv/6BwbAOOP394eGkm1170spzMlqbyoLJBg9ttnk
/ew+NIseeM1SeGesEzp2XRmRdlx1wPoUFcaPnhlp1S1QiYHfHb64+psaCyhTOGZVqo1bsO9C8THn
xAPs95Cc5Z/OfWR+wapQ8rtyxTPQFmhDpFSzvb7VQRmGQ9EYTAziudXnk67v8/KFeuq49iJSWg6n
sD8il6FMwOQnQc/BTrC9ZQBnRwiq3fhfiFO6It2qWUBAi7M5/lFQW5UjpqwydUoTkZ3WFN7Hqtbb
oaMzJzuosGNryIZBoIxUbSOfP8NHKyuRUamoOhxE6TYbvKa0bocY2q0xbic68Uh70Ld6HFfn0bEZ
q7djTKxSnMy+vJuRadYhxRnwfMcMLYaMgxh1trwsn/ZdUDJM5C3ShyT8Xo9BKn068RPJTeCx7hpC
xOeStDC+NmcLVZ6lS4JvLUbOHBYRtr07nOWwVOvNInc1XQ4R4o8Vvxt+kH6dceqMnM3SvWCYETYq
kEKIRfYmjTJb2eauoVxS9A/GXG62+vPKmvsjC/1/AAoq7KAxPJKEJKv0w+siL2LY7qof/aAAwJgs
mwdPLhnSPJKqA/AsCUDhVSdN8if/E60v1NdVGel/hxTNVDhNJ3/KeKtF7HpF+QrgBOEYRh95JB6u
nOdRjwZAi7jDOZehTDxvHcqY1AmNXAq10BqSS823Ime9bGObIHVG4cc72+P/Dk6zVH494gmKT9tW
6z0dRuVhglEqCG87qh7lkFyxxtKh6mHfk5RFpiBiO+dQ5JPg0ZX9lN0Te19VeDeIttWF0NkFZod6
Nb6Mysca1io+yH7c+6yVC7GkwMZWZ4ZrQr210caTR6Mepy+Rk9PZKg+sZUhedt977Zcp6XLpKpYk
3ANmXWYObCOwsnlvea083wx/mloK8I5+zoN78c/mnaDq+QGdOS1ARwOqy4hH5MopTgeXuhtZYgBc
xZY8RynALXwFqi4XyL3LLfdwcXW821xuUxOYWDxhnHMbQq6CBkgD3IBhYWhLPLQThOJt+maFcwg7
JfPW7rGctN2LChDQhgTaEcvZulonid3QBDYPbSxXNy3sHgxGvcm1dkZQSSo5rjQHT8EhU8WjdWyw
92Fbb5MgTwZETzT1z6p7Z70k8Qx3FLgdBzFjArPKJa/2JrbEEFGtVdQ9apZBJmA3tj2Ocl/7hZKe
kH0a5ljHPnMPeSSWfCag/0t66dnh+rjow/Jopv2zPzOMw4afrzSLlsrQUQFhqSS9rSBBQOJBJCeN
cdZShnF9TjtZp14i7g2YC25AZXYT6g62HkzhWVCllrRdra46m8hZDY57fqyAVhNVvL7VZ16mz5Y/
8BWHOImKZr/DPCRIy5x/LTo+kNBqRuDjxx84pOiO/Y5fppyJmvv6svc379UyL+k8JinD/ERApPQx
LKRE2pip08HBwwltpu3AbZ7kyO2P+D+ibN88ehuQ7avt0iEndtfYA5aCtdkVSG9th80U6Lv4HaBi
pdQ2G0bH+rcLFx/Rz3alwH9AGMj+mONm+rct4C0vzVOfAnrITmqzGt/HDo0rtycxIxnB4+IFuRjF
YasAZedtiSI0joL6rY69j8DpKarZBCDA5B08MyJfBkiruNFEA9JQbBESJdYtpNYsXq7ESBV7/t3N
YR7iNY3zWq0elcGA75NVyAxo90tJAjvB2L+2Q3T7fFpA1ZJasK+KhKENviF1SFTMdyGdsnG6FQT4
PgbWs958N7KwQ28DWYljPRJW19U1WyVen2q+aZrbc5CO22TtLIKlGv5on8oPKHZNLccRI09wypbG
v3Sq1mR/2zYZqHHXWmkbETRaBQfgAs/5Gtv8CUaGdyzgCdMwbf2S/wohFVvdp2N+VfNmBT2oxUBV
MqdYSR5kO95aLC8ebNewD6JhdfoGT/tIQJmAUBlz4mxxUXMRV6ZfjYE1id2LlXabgEWXdfw63vW8
vqxhpU6mCn7z0zSfRz0vRFJybFLIw3eVmMFEHlwkzAMVZyjndlwIRxDfAylZzVhXK2e1rLRqqAOp
QCxCuejvlosDn3BgGAagY5WlJ+T9cDDfflkb5L7LuRG5rhAHnFshKI5DfFYmHxXlFJgveswuUXgj
BW7pHdVstsy3fTDoOynNuMTGvY7qyaZdO589y9BLvj/TjJrNibxuEcOSdr8cX9UZxN2FfqppYjGI
+N/MtDO3LjjJjLKd1Md4Nr26SH2+NMxS1cq4b0rq0485H8L35F/FoeuOCZ+RDXs0laDi5Zn83/iH
bzIcUCkAuG4LnN5tS1DPUAdUnfBO77QX0iffQtvJ8Mm4uZg4h6cbKWLabPd4ImsY2Qmy6DiL307f
TYWl/B+Zx3ek6/Y6lM/djB6NcCOGK9MSXZCAzE8beYDvIxkMuOU3cc7cNZGq6UwM74TZMnBA1yB7
lIlxVf5c3YA7b4X1i1o5NSZZmoVQjBlcktE5JM6mLXPXQx22eEYqT6Wvz2eHDUQJeQeyRBW/FgnO
d84TwWVngkz0yiyY4ppYdg+ldTHEMnsVIN+/aEWITIv8Oz1YzvjqCfuxGKIZvEJ3fyDH/Q/6qEJe
wLdTAt7psK1mXL55AKsxzZ0iqMc3LyKplNrXYg7nCrjAj0XZhDmcp/k3oxZNxv1wRsUrVrXDSdpX
B7ncZcKaIRvhvssJistKdEsa9XeHmb9V436EFvdXa5dFZWJueRr4WWmePLBZEr5n5Z9qc7eq+m1p
Z3EQV7P+zdouygLxN+65KGd8P0j3mz358m9V+NmylcBZ/73YW/6zcxgzNQYWLtlPK2x9CfwJrZCf
GLSVpaoEaCoKNvgdahH8l3YqMKsBdJTEM5FetfJP5K9Vssyor6Usb55Qvpm80jA58K/dTEiOGfyr
EEM4fXORvXvS46hHuzQcbPo+cOyjISuHvB5fuZOmUjvBfcVWvOdHa1m1k1wysegRCq5+7q6E7fQh
Z8mKsAhXL+zwIBvBmrsuEFceue1v35Whp4Y0S4aQdZZsCPW08MuqZY7Nx5Cq4yIM34WVgEZN5KRk
yv03nKYoysvpZKg0HQslNrtQ7g/sWb8KJtxU0zO9pb4EwbXhUssZBc5cbv2VyDdZdNX9l6IgZjXN
mOw8Y8Zs1Nb/ZAmNm7X62XAzKcW1TDK4ROWgRiqVzX6QgCR+rT1rOb1qNMuZTZkHZskhwdJgFeiT
sYkGCuXajDql6iCLQZf1Ls5e32WmpLBEAxIu+7LKK4Ji3Y6aix17e8nqKHqGNPb87e3pzBRruh3S
j0WY13CcvkJDV63e6hntNsqq8MJNtPvIDXNEwqOCqRTILdRcNuRN8bA8XRhI2J2/JiPQmeemVs1R
tv4c2HukqFbQP9beyLevZieDCNAouKOic3xfvBFuwSkIMYb7/Xe0YC6In7340E3UUHgx90L3oI00
kZKilmSztpNhybGsFGYYkc97PTlbMnl7Qd/Om28auS8fbeUJMOhkdL+hWhD86lu1DKt3l5i65SGd
0cJmRGL+ladB8dn+KXnl8i+xBcwkE0Njtev5cjDL67POYDYdtKxCRGzVVk5DNQEvU+8ylsMPsY+L
8I23TgHBHNcKK7HTQd0iyzjmyfrDLnhhGdsGZ+YeCw0LOG9tlik6i9wXyfkVfu5nSH9X8IupMCFC
Pk6Lwh8JPylJp4mRGF0WFFhxCPi7sGPVcvdWmG0Ws6XvgzTRWvQu8YdgbPsnOvnOp7aI9hQQRCZs
mPe5gxweeTg6UE0yT+fx3MnRLD4wRpi1QjNUvPl6VC6OtjRmUf0vHWjwyVQRUgWaUp+ax1x8ULT5
jZrHcueUrBA86L4NXpIPI+7Ya01VSxkNfesK0Y8euP0UcjfqUvhoksbdp/ibG/CjLACDsTeQSnrf
ZaA6t8x8OBlrDPzw8uZDQQ31oQOpa1I3VD67oYP7+/hmNmjWY/xFu5+4IRKyDASRJVQHSvkU2LfH
GiZshKtESIiJumRwYJK+TpTJRNafgfmM5tsA9X5EM6iL2G1mqnUFePLS7UMj3C76bOlNqQ9r+hSe
6YPS6ZNEULJUTSM4LyZKZcWd5KS+BfSc85+jj2OdizqNh5iQhlRvr7cjeSyncbAcLfC3woOXG/gt
3YW/t2kQn8X87gvhn7/M67nYrRWw1eCuL4uF8fNNv1VP+IV8i4IlpmW2LJWxdmN97/Lc+qJADx9J
++AWiUfxxMJvLSfqfwbt3v3sMmDZX/6tiaFubobYkFzEN89h6gEq/dHS2+8Y5+StTnylKR8yFj/5
snT8mvqWB/WD0yh+1/eTs6iXbWK20Ad8A2aEDnG9ijtOH+APfG9x+4OdPB7uwoos7aisxDsnp2Us
TASgs3hElnVVKN8axtrFTb0jqi3sjO5PI/vx1NM/Q7Of5XKhqr2l1CvahTILf7q5QfI4Pm/dsfFd
C//oVLU4TnZ/rWkOJFNLn9ePzq6xfckSnQXX6PeKr8yfAFpwp8Nw3C8G8wG3uHRAxDoUwL4mEJOj
nwzE4w3gssMh/4NpyziqBxyau7+zatFQUNokSOo8QBdJCWEc8JHcw+VOCa97NwRDy2ZUuNucPzrp
wGQFJvR5iTFgARvNZQxg4hs9NFUkMt/n4cHRx07CGV8Tzw4jk7v2lOCU1tERxYZaEPRw7NsCEs28
wB9abu1+xWZ3/fPCLp8AbzGHJn5JlBTEMplN5EPgJ05sz0TPyL3K7JU+aALG4mnnF11oakTy/ADn
0DC0+xk3RrNwa8G3XKCAZNpkxaXAK7StTiDZ3uQFab8+UzRnXUTDyqIRut2t9mqR8QCUa/+rAx2Q
o6W8SgWjdKgo4tabauS/kPW2eDYWPQvxBZAE+sX+tLPZSJVlWt78o6+WItqg9GDAzmgjgfp1FFqn
P874G8JAk9dyFYOxwCDUnZeEwkLRiQ4lTx46lxLLQRWzcEdnFaGaLd+kWloJL3ayDMMEBmBrMX8z
BUdgm4y/iILb35yzJAEeLtA+SFpSppE06KH+RSSHKm/7d5YzE1nco0mPaOXxq300/3TXV2CCkmTy
HGeY6KtMuYQbi0KtHotmC2zi/Q9JTiAfhG9OP0AI2V2f2BwLRCSl4BYRku0nCeIyAw8Q4SLUsjl1
wEoPYtlZKWfEZOUffkPnLdEKB4qj43GUKDvdrDHU7sRzVkqmICYV8v0H7UrYKW96iNswraBnfbHN
CFk0tFbfIVKofY0+6+B0/tTTca4+jv25fqED16vxyVN9NMsomcx3orglqOO8tOXw++019kwVmWTQ
oi9N9EB+GfJT05gDr9pRJVxNM6MTOwXRaRZNXlk+36Q2/FIuM0dZ41OF4NXfAOQJEqXVwWbInp+P
rgDcwPaGcsHs0V3MmktpQaYnF2s82X467sCeTpDaJ6E/TOkvNNRdifSnK0BLKN2l+jFfATrcZPcz
MZePDU4N58L8KRwNHEiNkhxNTUFXvIXD+nw0OgVorG6DVnnNjTifudbjyWf1s99rIOYURv4miRH/
p3whpvRSmil7aWtCLT0zRSIYH/RH079lh1Se73Ntr9vOhN4x2okbm8v78U6FwIOPMHyQn5Nxltvg
4i2vfOPnQllA1a43Kci6/1jRtRV/0TpU33nXKs0fgrWJEbq8+dv5Eu87dnL+suo4lPVrC2hbB857
kIiHuSYLpX2ih4XeBiEkfWLpCGLrvLk9seaTFcb8Rt/9EOalCPnpWJvUrobBIQDJq/cIyDcy/2yJ
2xBKkzE2FOOiqfF1DpLwsv24SzQVQZGKCAHGiYsandSk2JxWvYf61HnrEwgE49wH9bvo0CsRWDJA
OeA+E1X8fH2HrJcG101aUBY3gyLdD5I77mjx2xOxDqgVMb/mwE66CNNh+9VUXJfB3YYbXZ7wfajy
joNi3ifTN2wOkvQLnOpq+BY7qX3L/RkX8A4j/ScJPlyOW22EVt6q6CJUIIw7b+4Fuy0CVzSFYoT0
L/5PPPbQr93ecPCJ0JNpu7yLHeAWhKL+XlnDU0y/3TcFiHKycbtrEg9zg+xHvt7+nCdOczk03Sta
66fc7tW7Am9kAP3OfAR2FM+pAXsSqzSJY0ZTBLmoe6bL4G6pKLaY7mm4FqnKDz//g2JWibam+1WY
5nIfsPr297uY9d0iMUIxo2dkrQNIxVNptUuUKTy55dwVnY7OIPCw6I2rhiwnT+DHX1Um2FPvD3+a
U/Wcb1DOYa+bDBqilIaoEKOy7x2qHCuS6+FKYtNR5Yw7c1KuwaSxoLstdhxdFyMQe8G9Iwar11w9
qC2tq8Fj+NUVvmfjEfGaMmJeNBtNF4+alPX3qMFUiDaR2Ft1RlEBlxfNCH8CWvuUrtgcZFn6hvVv
RVKi9E2I2QO8OiFxfhbfzuKJp/VhyeJp8vqasqgZjcGNCwuEuRFADIihIx1Yar5mNCFjMo6dl0XF
8Jv5Pk89S+okhiz8XElGM1xe++dlR8pfmKVwvUC7sdV6cskWC9yYqu6SyhreE3P5v+6f7xvRW7oD
hi8beDHxeUtwbdftO0rJmht3ODnbV9JWTVfTH9fuhtPqgdj5nYKR8OxbcLmXQVEtnNaMIGzBkN00
HNNytCvHnLY/6bzQ8XjvUw4MPlHfIyH4NSo9Sm7BiAkBJ1bPXzsSuLYshcr+W39pioymyzZLT8oQ
TWCNYzAsl0LJ0xCJORT4hu9oeSHqnscIFIxnU+WJ6wN1clwo/UTqymC4hTPEIxm7DajpRQaO59ZQ
rd44vTHcFy9SMT/6o2fNd6VU/U8u4STSB2qnxi1OQHDvfGyjsa6hrlkUhsleBycrRXjVl7dtQJ5W
nJ/RxhbtrGBmRnp7ya8rC22RS9A4UlR+E9hfWOICaczymEkAJGbi16kzJTgpEESq48zpVKYoDu1L
u3kQ5X176TO+GZpJUnRbhsnUjbxsQKgtd/WAAeQ/XCIHwtVAkH+ewXAzr3V55tDlAUy5Te198d4W
f0vfoaifZA7Pr6nRzFnr426eURqQSJIPOFh36paAXXL0SI9BbIvdOFgYhQEQtNjYdERiRvgmlKtv
IjLWZKjAK8gHz5IPb6UIhdQezpUuif5Y5c0FRGtsxkigI684U+FBybOfOsGGL6DgEtp6Q3+HEQK2
VvIsyUW09UroZgaq36LiPjnLXYUs7ID9AxKqRIuxR4mAodxu2sr4INKexV4ezofNJAxvx7Mo4wKh
EL+nOjrMHQe1mquJmf8HpA0ki9Vu0NsKK3/4P68pcchjsii2WZaodCnNKnwlWAnlo4ZLYBePfh8i
g4X5e1GBcCb2e/dI+91mppV6SMrVn/all2LyfTi0x0V1W11QHwCydsoe5/v34BNMX8us1o1ooyOB
5Hrt+LFH0hNN9SntW1N31rWHCpGC5MI3ZoR5kLbnQNQKbHihESnVga8LvZmexEozy5jjjilo1Rqa
ErfbWNeXGzyjxGquOEgQH92SPHsvzfAZ+2T67UA0VGUXN4SUvOiW/WD2zl0hZQf4Za2ZaIrlGsQK
49uZb22lslGtFgjsDSvwWzhNSSFqIua4kehmknlJUcyRzNmE1CSMc3RhrPf/6qEUD/KtZkDbQWCN
2yiA/ty07ACWO/ZxaPk6y6uwOh5f7rQlNC/Hxu2UOQvi05qjOisPmmrskesPljaf6u9qHmY4Rimc
d/BYmj+IQ4296elLRSa3GmF2NTjkcQHyOE25frtyGONYhhXP4+u0xoOO1IIbkc9pehyULWSg27h2
zbDFHQ1tGQ/sP52OZjOj8O27eF5qF8NjMF/QexSSCYxMAZ8vELU51xisIShCJ8RDRGsqeU2x0p1h
S1xgzUb4rBoh0HD8rUjn88z2yRV2XDMg8ABSEom+UbLVmfrT9RhJp6XmE/8F9HH5fVeNCc6oabHI
R3H9HAqDVY1m/j2hKqlVTpTiPfIBWQCLXxzFd3WwQtRyw/cUqa8s+LrGZBBlJwi8dGHvt4YpaNhP
67qCff6PfvlfbWC1H7jd+6zvGutwmowsE1AkKebzuDt1PMGkqSp7mjGUy0WLTeQWbU1SPbPwKJai
Ma39qYkiGNhm99diiUyCmHn6/DzJWuLGrcQH3Lt9W+vr/vKanoaEtQNFAJlmlczcVHXTIDKOxb0y
HsewPsWlUe37gG8h1au0V5g7KAIkCmHvI4XkyRQff5tCAJJ0oL9b238U6ycGdl2BO/hSfzfCirP6
3bdpb9sGdQjbuAJO+ZkGsOXW6P26oaADJ0fQZXTTBtMvH01a/ida2jPG2D9Xd/VrgYoFRdgNOKbg
Az0vWDla/b172eWX6wLcHuxCZYTHna93M0Fyu+td4zsz0qa/yODZv7OX7FNJhXccv5/Q0MLvAIrJ
9qmGl1iifHompbd6ZLBY4LvlFvJxnYgn575nCEH3KyNGgTCfRzyFSs44oFC/g2QoUefarhybU4Wy
wDSYIt7YKa7TmvW3wIMKvAKVj9MPKgVYnBGcCiWLnQ1z0QqsjRJWJ413zlNw2mFFAxgr++oATbrc
iR73d1LDs7Cb2yg/vwdU3Fq3JWlkod+OBy2hQQdqTmaOX8cQ6IxGLBwbhmIumN0z/eWFs7FNxCQy
ItjqphioWR56SU3Ta+p5yropUKu/LcXR7G3XGnC9uBcRVDbk3uY2MFRm9P6fkE13IRqUS1TAh8KO
yiJRuJQhbrwiStE5Ym1k1vaS/Z56DPItcQKoZDkbhk3dKNtzjcOmpUJ0GdoMk+sdQkYhQ6Ujq2q/
K7It/R9ySNiDpu7WprWLeMVs/JE5nPoTQP42pjgNf8HTYmDVJk7exRpJ7rfEroxyEU5zXjAu0+B4
8cyfShwcgddGEr+k2EBRLpf/cgK+Ead1o74MHhfyvSTt51vaWfmITRTa1nSN9DBJ282a3MZBYMgx
tn/LTKPx4WZIbqWogVT5Qccs9cb95KEYUu8ivfWkWEydETeYuENImlrVJGIHszZACSe0wTtxAiwD
B/AkYN0W+kYkGU3jjr2xuWRTB/8dWr9TvjznObH4GwfsUk/MvpI7rqPFBzBhD561Tmn+lSn6dTYA
opZ4v66J65qQ5sTmUZTJ8FzKKkrUPLrNoVSxxh+/iq69hWGdVlaK5+pF4HMniKzRGDRRogjalCIs
23JWYMN0JPOkVF7BZzyyVnmWDrJJ+ntWCBDzRJFyRyEK/jqliv0ZvNpQ3yDGPESIVx/Fj1bK5V5R
lz7ZvmmbW7I05p/JysJdQq9v15XL1QPvYwiesH1j9An4/n6TlMWNHFpx6vLmqarvkzdEUfeYFtnZ
lNMD+MWReq04UDYTVRAIVLPn6TvIwdcNp0JOWQqBlcr1LXoqTIPC7zB1u9wNKz4IK3cMrSakgJmY
gj1ui0G+iqFOJafZA95s2R31Kb0yeBmPd7r+1uQ9UuAhOqGmXXnChqFnHlIbnuTDmNHBiOdnW11F
2BHURyQ6k8i+FKooRUc2IQGQgTzjC65ePI3IHVLOUmRYqOgHuC5g/clKQTRq2X4tsAarJRr8/H8g
jdVAfRLmMwlBdtFpsBs2gJvgyNTQ4MRjzE+G50EHmHlPgYBLPojrlMk5Gs7wTm9wI9D47OJlCcJK
gIcRW0aZeUASfPX2g3FCxphAUxewa/D/HthfKkJuX0cMyRHmznThdUua7KK1GaqxHSfBgC0t5klv
cqHIt0c1ksqwkgiArxv+zS2LdLgKQEuE+xDLYW6MLgGzpUHarwD9PnsdLD25f89Cadh4sjXF7q7+
hrQUG2G89F9bLECZFKKcxAAw8AuCnixE5rpKNa9O8P4Q5W8rI9F5g4xbM66SzVftZS2vZHAlD+vP
gOdNuCj6eEVkytIBC44FFxY/iElAyqLkQbILf1Dh7tNDS5PaRESA5Z0XGRW9Yf9Xod+txl22Frvf
fLHN2fSIqyVGqSqQAJCSkpT2D6Zhmr1INnKEjhLc97dYLWlOSuv3jwQfrjAL+F/JoTkSiWM3k7xp
ljeU9l63+YIm0MaUvA3hSIvMl4yYXUnwkQL9iRjMROilgguMuyn/Fz0iVPYOsquyPd6wnbHi3WAg
IskiJfruNzdAl5gytalGE7fgCUKy0xh3XO7uleFL7dc8D92LuVTrMo1adZ3bEeKRmUevf5n9g+kc
daKvmOxxby9wE0pZJ4YkpuKtweiYSQ1iABrZgPwBhGHKIOSs4sL1YsmjXMehYfxYHnv5RadqREVa
fHnrqIMUURZMy/0wYrulb5H3nSjUnBcgQUhodXOrWHf+NJ4m5G114B9sldXcOxy4xKCpH4rzlrsX
3xxwm1CvVnJ3lo/kPJcicm0KeJtz8oNAOtZIxI1jf6nMrPxvFC6cUWbw38fsAWi5u5duI9UzjGw3
f+qkelsMMUt9oHfBnZ2vOlVgSbqe3yYSr6ACw4OMcPVeVhrgFO+uMvyHpzOW4Quo8DNminjx4gkv
9qFz5tMC4C3K642Jo3xcJ8r66YZagHAXVbVLUJ5cHvNXZOChrcbEgZFXhFMWYLoB1+rvmWjIy49P
advRZ1Ui5derUBz/L1GDIfa9GeyzLpkmCCc0vfzIvqIrI21WDIpm3uGe2AVpF6kA96Cnp8lSMNpn
W13uTCk/cvtPRNSkiHo5Yk9CKDi2gFboAC5kWy4BzpDCuNBWonbSN6zclHbIYVx0sXcqD1NCSUQ0
fdO7ZcTzF5jGF1n7/ANKqG9FbxLFvQmm4bDjk5/AsFlnDxYY4woKXcr+3WmwqaZ5+FOyIpwRqnm3
8X4HHKh7BPo7e5yha6NIto4oEiwY0sRytyIeY3HXL1TC6vEAMj6RleLuikMfNxwO2WSxB6YnYuG6
ZQWYE+cW8TvNIKVjmOCKVZVNjFNZorMObo2RA9i6iSY7hvM+1H8AZ8msqgafFS2BoOS2fOtfXkX+
DH+JMmkr3JWTDhoOwN+tWFsh3CmxMUzbRduFrjUdNNKqIHtuVXFmYE9VNx2zT9zg3rLn1xrHYEZE
vmMF8JV14YJtK5jPEyil7CV0n7Yw45ubHVvXl6PwlLtvffYts/loijvgXGIXq9lHy3X9Jr6Q+Xx8
DasSyceUdzMUpC/S6UB6qM3I99j50RnwGEiIr74hLp/kKh4lcq3FOIzl4vfywNMN80TjpLtGEbrN
Z75q0k5KkHipbelPuqIPniLrK/NT6vpQX0+eQxELvCTGYQ+255vsu6edw+v+XnOHMrW+6Ew9G9Sm
teCe6WrHmCVBK+4LbQjidB7x3BBvGdy7QaApOtAOy440R8b5vTkh0uOfUnnj/KhbFIqdFe6Ta0QX
yPuDe607UVQKTGXburqgUmvqEFrrTFDLVL4kR1PgLeG1+tVVD4D1RmmnnCxqowzfP7dGTZhDMRgX
tOVdUlHQwtIkpBgDVkxhfWIJsnM0g88gnGUyZOIJS/68Z1V0oF3ovd+tkWMTYlxa6FhREcu1K+mE
jHv53PIuXJWOhxXae6nHYtbYJhbFDuZfE7RsxFGHm9v9N3EMhyBI37D6ZR9HPFa/nkBRXhYajmP+
bpea9WO5tlrnFfUruIy3saFC5xWJIJjXgMrdwtbToZm02rWp80MWBPrvckSS1dcnv27MwT5yMne3
QT0jHUkjC3d0hT8MTMaCm8u8Yxt80JuJE6gfO8a9ui/Acu4g8WKUS+24vOTgstD6UftiFe/Ss8PA
f20dis7AzZN0HRdiSgyxbtg/51HbSz75XYuCexfiLheoDBAzliK8GiALyjYrQW01UPc8PxRpx+Gl
VlR9jETAR4wCoHmd5QcgnMaKxMiR2jfMVqUzhUOJ7LDRwAjxpu/dUe1X3+sIcYpeFc7DSF6zqCux
IAhD2DSUJwjXT6jgWcj09CDi/6Krl2AMeVD4Wye1b315h5xJTXmoJ78jaBK8nwSZ+BREpJZzDtSN
CQ8yIrvT+hYUmXcAUcz4w/cQQ3Cl3046/awwhLgeXlEjRivMkLy0DcXk/acWESG5Q5uExVWcpsfJ
1jpQ8nqisAlcPCASuVUVHfaYKNAZnuyp4bwWOlWaAqWqQHEnHobhvjh8KfQ64ztNZaGu6fEsPtl2
jrj6yZMpQHWayjDNbzkx8Re9EgdBT0sOQ1g6Cs5E+d5pYwjEkhrrYpWsmlUTVIIAxYVjmoCdxN+d
IMLV9dC4C4FwnLXsxcHsxFAqSn8PFndqOcEUCom90LYbtsyJ97+FQLtUuTUk8rxRqwjl7TROnkmD
LMguGH8TcWjOMIoCRdwxWbDxS8PZ4+FBe0mikQzWK2hafh54hDIR8pPmPSDfv+/LuSJLRfSqAgcs
ixWpYpi9tVraGOLNpsG5ZhBmLkTrIfWYdSZgHFWzfNUAs18Gp8berqiJDKRb5IKwnzboHXisTdfG
+8oYkbwjKYwpTH//P9IOwI8bPEI/wS+eHXmjtX4Ie2ddhW1BzpzYbWnKSPZ+07CIVCmln7W77fgn
jF3zFpY+1+jTX0GusB8ClHmtwwOc8tdrGzxdg85fw8yiVla3Ofl+7eGOfvdTsYfwJXO6rRpsqd6N
op3U1Auz4PW809A8idkUf7DiDFGUYmWrPOUhnNbdqk2IiPCgO6ARIWZ8k9ZZi8o/PsyMUK8iXGC/
UppDSJlSKyeK5c1GCdBupl3wFJ2QPFQgXz7P/SmxzONYUV1D3akm9zgkXSlwU2SF0vi5YtGaHC57
OCDqW0vasvPAiERzsl+K76LQM24bgT4QB7I6hyM/lf5fTkTUo4FyprLNltAb7vt++UR3zm3P2ng+
tt2aReLStPtZhs8CB5D398nyqP/VMDSUjWFTzcPZsVZvxT1jwYveAE8JcZLtLIICywBOFomJ+EvQ
XGfAxs7KLsYkJPnGcIF0edJo/1cqNKiscu5ArnBYlpbJOumWlg8Iqh8z4w+5mDWtuzlx1pdw6dyt
0A+rAnA0OcjQKc+DYn7Ndoj2+MuI+ZXWzo1w1siRfZ1nlpK+R/OTqaH1drs9QOsliQgsgDzVxR3q
9VsoW3SkPRlbiMt3ntewJ6TmWlPjHage8sM6ZcfwzqRohA3ElCgIF+jAEb9POg1mDPLYQ3usHhnY
xH+JCDV2pKvrzNOWuYDwAP6+Rl53xqWV7H0w6iUOKjc5QfvjGcuCwuDRRUbbI4HrdQMUJAJI2Aue
gvHE6AvO+tufJnzVpfYXuV3JEWuEKU+D0Hwoasm1cC36CX9pu3eKzPBEzXwD6D9QrR6rmDAUDGFM
bsT8ZEzapDmaUl4S6MapLQxOk7VeZYIV6AdTfmsTUvvXLaRTWWdXs6hXgooIAJTdWR6HvTkhi44n
uxEvkSnzhruxkGDZUI3GZjQ4hi18aDXjWH5P+AvOinaC/fJlOIVyQbyvDwvuwoAl1DmkZMwCLr6y
amvGDIV1cfKbH+pbK+bxMr5kVLLjWNK8B/HrM7CtyL4gFtljfEhs/7e+RdI0bnTSPpSr9M1dRQSe
mfDTZXx7ymch0HEFPrC8KReDNW7++WIZ2gFHpvCIWfcm5E1t03qv9legBUYafBg9+j7qQgi5+god
NdTVaU/UWvvW4SWE49hYCSkTREkUk57JWVN/Eu4YydKR5s7Zpk6p1oMix16DB5s743aioT72kzkn
72mhq6oBFU8+e/HNJtWiJQ08YbjrtqGy704P/1xV7a4MukLYmhpkrbvB7UKMvQMZbBca5bm+TfLq
xk7gMBOabcneZrYyGwsbScZsrISjMFFdslNa5Xe8sadKDv7SKfyRHmYz9FPtdSB1GqXylS6YJiR+
WtfBpMc+3vCJnyAwiw+ScFA7DmrLI0qagzQA/U2GnDsGyIIZvYbASK20/RJQbU4MogGzPQs5fWl1
2oGjDXa4B0k4F8mii4yuTICYpVFtC3WeCmi48QSNomlAoPYaIj035Bw5EubAa6oudLUFQG0PNmZy
gGm69HAWGAT79qYWEa5Nu+CGE7iXAtM7IUZkJWrdsi38nrzbjJtMGj2sjHpUaO69rtDkcpWNhJ5Q
TDT1Bf3p0n+o/q4YbFzl+4PR1i3EFpIkgNqwU4XHy4RxhzpVwyHiRfYrsFijbgUfmHyCAff8NclH
7F3IQ8hXno726vZwoTtV3hnNelL6mmBE0Q1KyvV+vO8HiqjkEBe5BJSZs5baRyxCAom5Wyit+DhX
sJK836hy5Xftw3yLDa/+yJeDCK5RH8b4YDNpM8Ah0d6TZ4FQIi+AUvk72O/xW14Agx67fmAaCKl/
YMLYN2AwAeiWoqDBZT9lF57dOsp1ieM4pLc1eUcdwVqthdwmJf0xvnejFgiFHNzIkuh/+rDenW64
pZMVq09UaqSK2u8RxjWvpdF5Y87j74NluaskJzS8eRIaq4/Ymbz14tF2XKaar6j75vdttn1zRIS8
2PbtUXppVO8v30F8kXBbX1iivwGnhCZfLFkNQEfifPQ3kuj9hTU1F+HgtoKLv6I3AREjXKOVWU6s
LPzSaWXKbazonpytDK4ugFlBhjdxEcmkcbH/eu9lanLSuRk+BVIgTmEvwY+cQ/9BVyvwzUuLquou
Rih53FyF/alw6w5nP7HPNXq2ZhjY9qc9Hr3AVUsntMy+Hmt0WqsIwBU00pazICQF3ejfjsR3sofU
fpNCCeYcO8O+Qzsi2uvca32Ydx9ZTks4z1pSr75Lfk2/CuQNC8znANanG9zhmy6fC3TbFQDWE+Gg
WLVBT7xx6h8XJM2Phb0H4kTK1FNPfAQ7T7onbdaKKSiFauVk2ASnsCaVGH8Ma5bcsG9Q8vRzuRq4
M6S7pWClExEMnkp5vvBDn13Z+31zlB/FyqhWCz4m9+e/cZHfkNh881tYHPEwaunHxK5FGF1tmuk3
qLY2hYAoQpl53rNOftNcXlJti6sdH8SMxBME7G8UQupC48wJts/Cqgey+Irg5jPjtsSgyx79Kthb
XadVAT+E7a7vCZnIToljnzlZSDjyDO/o0/fXi7uwAsgfIyi2G2u3813C4J5JqU9x6rib15tSZPjU
h3DUA/WbGfZx89DgZwVYpVLtNmOeBC6TgmdUeGD0u4wBuBV09SYvE+uS9yDqFPm0TSghaZzoTGiP
GLtHZpmbGwoyuKQewCkKyD1NF9Icw91QbAFl28/HFs7k4F3bcOAvxlG57Z8eZk0X0Cc1M4YkKb8G
sZgo+VfKngxkHY9rRZTJpA1kC2d6fLhDjTMVR9kg1T0SKOXq7CSqNBaX6E6xlETkVZ44SEKD7/cI
dfZv3puQdxQ/mMn5nD729bg1TciQQOoJvFQapFeYRvcr6c0WRW1KilRJnYebvVbLn1bFWI5YYd0A
nHygNwUG2/9X0mBI9y4lNGpNqiE+xq/14ZODh7O//aezLR47W72FSExxUYynSknqrvaOSkH6Wqgw
0e1XE3ItEaV7L5AYRTQGr5XqP5MYtckxPMRFN9MrWsY02kTpo9lKSzWT5eIw1aziQ+liIy8OqIwp
u3ij4LnrrB/9zcXR0l8XWqTEm2dLzE5ue+JhoLcJjNJLgj56iCOD7ILQTUJccWjMcMsib3Gl1TGO
6ODQgrzPRbxTkbN0+nonTfYYgHUlLdMx4qu1QyNsLu02tiJY6WlBdc3QAG+87/x3GUSRa/5f2D9B
Lmvu1tt8VAgdy0PyT8eqKRab0OZghTZO3kDa5gAw7/AY6+snsGHWbJ/xQFHrmcjcw6/yp0QNjpB+
QXaZRmyHVxcbu8Qy7cIJQ2dgoWGsfj7f21/UqqIAsuY8d7nB5AsQAB5IK1WSwx+mxZlZXI0kytU5
TN9JK/Ov/0ozIlFH2veFqngQHCnCLx463OiNf/WFsnbcFrvxC0MTZNHvvm3TYJ2c5LpB+mHeeP0H
6P6nkUt9CEFHUkczD+55MQxilsUNVT7stQoNlVAysTfnVF5nUY0FCj552S9d3T3bAHD61kQNdt4y
MrjZ3gmeUxE5zxx3s4vRY1XctEaja0DRj5MzfZ82sd+XAGJMdmjHcfNP5hp8U7Kggj++KG7hr4KZ
RF1KWvo0hLZplmDnsAFiGgBEiyxmq+ZsqJyovDRbzTJCXeK5qcVsXsKYR9YghvByo5j30rWbUtKe
1wdww9Z4AAgltyHYMwpsne8MgS0yizac74CUoYRVbAKDdRyAdmHl638QRI40T61WO1AnzzDekUVQ
l2DxYVKX7ooTSqASYdEmiD0vj0k28vg0QRim1AA/Oczm91kPGvKtdmhIN9bOxi2mVi95TB1V68fo
Viz00eyVH+6IyaCCYOf+WHkqHcqfePuEsztfv6UJJMlmme5jcaiB81aJ/7Ynn1S2wDlIvioODBs3
net1UQy7HwpL9uGfUIGt/CDIeter2KoPyXiekGk/6lRS0WZYsYacuWBUbJesjU3GiuW5WXQSSo1E
WLpmvw+Lk2ZRvMn4p/JPnFEqcYVCUfcW0GsAS6jPceRCcbTOPlx0gPQe4mysniYpcvKcOUlfit8Q
dnnv1mPVi4bTho5pr5y+Q5CZsLXEBxdGMW9FpnTbbEkm/antsfFAVZYgwcPWzqLo91nupx2N/RM+
itKkUik8dEw+n/YH29pt/6MVlV5yEJalc2kAE1MHFghC//IhgLnQoSq72PhhVyqGDDmuJ3HOTklI
fKdTjOSJp0A53Lyh223Ix9YvhVPR/Vsl1v4hw3Hyi11KbyVN3JqWpMB0OyQe2q4AIGfu6JLy/aYm
GjHQllxzg1b0B6GQCAOQlixPjuByrf1IqTFA+n9HcuUrSgmEeRsuPo78DMtb+0iHtkzuUu6r9aSy
CEXlpO2KGlxCfd18A9nuzOuEvA8woniZlEMt2XT/haaI+mx4tzKwi8sHrbEu94TcAaoTnVAWFxX7
aBtYy9eAOU7oCjwPQCRI0JFnCVhq7Tpw8+6m+wvNVNibCDP4vuvxDR6Sf79EbWrMQTidpkfUsOtY
ay6pcqucTxxsiOukz0ygwdAzutYmHsT1KiiBwA5NNVdaFrMzlDlxddbBiOTZbONv23S27uy4ujTB
gGXTnYBsILPlYeyuYSOqnwgBUWyPC0dSqVD/7UM0IwIF0rUsF0MGabq+kZSyD5wzgCP4upERldNc
o0W981hAH5nRPRDp8vrwSTDo+GrkLudN7aAjkvYejnqWs/BTdsdfAzmyD6f8RY6TVuTuXd4oC6sH
UjK6v/QKGcBN1s4oP89r01ni/XoPtwgg7Dbzm4ecy9Q0Tx8q1Wj0fyKM0Do8GFDXGAXKL7pYEZXC
LOjgYb3wZ9CkNQ9Msoyo2myUprUKzA1yH94P2ZjnM0RJKoXateO3zD8hdm4eGOPVAeDgjutIBFIx
4gE+bHN51gbsG0+yfrkA44OYqIR+lKytswMfgdCV67+EB3MkKSjhDSYwZIc2VtvsxTeQHTmHB5to
FWTbgAagK4USXUwZl29Kd+7Y6joN5XBI0+AsRhkDGjpLrhKgz0Jzz+sxQz5eprsaV2OJzahIF/D9
fH07O2ZvXSYqOxniXD48+I+KiNIWEJLkYgdub+jBsQK0w1eTrG9EhSygDJ3KsvPN8Pb/GpfPPEol
ztb7MCkfs3lo+gSi1hzIcN7L5uJvkdVHoPliQi0IMjgFomEJhiqqBJ/EURsRkYjKT+rQ/RiIekc4
TaByhW6oNBzFlulmQnjWyeUXIX04KJjlOClXKw4Nv3VCU4z0ltOOo8BFYFrh0osnvN+iQ3hTpK0y
kOtpWwbOzNZQQHByLSO10HhB/7Hq0KVLrxRbLKl17ZxbkEZeWwbME5quyktC9KYmDbUcLbBv7lSC
CZVuUEPRdW6vFmT63uiB5sDS49TGDFLKAn9wzmFmEwYPqijPQkrUY/CtkRh+coJP6QAtLjKz9f5P
yRsV2T04TaEPQ+LmOUppPqMihBs7bv5XJJep6v36R9CxzlG4NlSYMexxbCKqNTbmu296LTcsnj5b
zCgEg85fSVSNcxpq5QS+K6PD2YOM3FfR1YjDUBhkIXmqgbLDp+0W/PQYLJhTzt92iMfIPVcs4jjN
wfkswDDFkE2cLkCkAlr1i1MUxoGCKREXqwF6xP5Fpx4dIXk0KCcyah/bvW3A0Lb46LhCu5ozMDgq
m2rXfotoV5c+PrXzhe3jdExu27uRLV4cYbPHtSEBZJ1H9TWU/ccis7UZsKGtF6Rww2zNfOHXZkpX
cu5ZbF5lLgtuvU+8SRhfXB7ySrV9hNmNdqhHGKHSILBmABnWXCuG5u6Fknsb6PfTA+neDPfrDA89
+3UqYK7D4+wKjafDQnihdNnGiSEEwLErP9jkHCcIjSV35J4GgV1GoC4/yKwQwVtk8/tYq1A0j9ae
Fk+1tnF/Ps6FDfwKmrCH7e1BtetM7zqjszZKLnsZYxaFZMMiK7cqmBIs1v8b8DmQomQ0a5/yarUM
jaEFx+ZWA15bgVjDoLBZ3F5TzTet0bUlIcH45yo0qcuWmh9lUiSZEYksNdTko4lrvdBDrxAqx1Gw
moBfgRrXWGOKCv6O+1wpOhB/9HQ/m44c76xrleIue8d2pgVruGJ6xx5EIenKzp8H28uvbZbpHU8D
KdEWscUq8fobezEEqRVkmR89V5lD0/ik96TMIx8vjxMBvIcIq6PjhtGeU8LVopCqfWSM83dgGtOi
mipXDK+2iFHIkxY3xEaR7aMMQTFfSILhlPZYyTjuiZGLAQ9s+NJDr9xkzzlp5dnBoiltCDbOfONO
tZaJ1RoDF8595D9BZkrGIEhibnVyIj9JvdMDIxill6yQR6cpLP3fGyWQPZpTYmDlgKX+Egk97xbK
FaNYWja9b52kirOhWcCae4feQtiGyQm0OgijBS25GdOpFG+4tVjR4mrtdmSxNz2vu+yHiNWgyGuW
WAc171QLMkj3DRXO1SLK+rtzysIwqAxaaPZfLdXJrHbJyUeydhTU4cwFfO5xWZsTv88tBczihy56
YDehO2i4xfghbUxpveuf4ZEbWpSSkatt23fI8hzASFQeKl+YRTfbGvXU6esEl2bvWY4ytfTN5WPq
ciPHW05rU3gV4527cAp2u+86IO8mYHmfVkJOR0RCX860ZGQXT9+f+dXy75FFgryE5xWnNxwxE9e9
Jiu3Ac+8ZhUklok0Mjc1hJa/v2V7T2/m63s9uf3b1tpqqdJpNXfJOLflOg5XYOnyzEGjYyFE6Hgt
X3CFeZHOHe8XD3RfAuzor6BSfpPpe1ihTjYtEjL74GHZD4tIob40Lliy1Jl9ykotVZKshaU36JCr
cKc+gC0XIsyw++EvzyGDclSbxx6q+ftyiQsrCvb+AZCBlucBIxCFsGNmpN0NxyJJoro6RfYGnGhq
FlnCnGoSsrb2SPjsK8BZO1CXQSJBumhkHzfgaNQrm3rTezVU0jAAwBeBOrxKj1VMjUYx8j6l6cNN
d1Wfqi6u7xbeTGblcXfOg0y1p4kzxiF/zZ+PZMm6su8rXgnvPqfvI2pgOQnRStCJkR+HtIDmw3wP
f8fbEXkI6h3CIu+1Q7eMJmbBz/zDI69wEU3MG1MMBIGbXsANcic3NNgJS6jJA+izdRX0OJmDIiH1
INxSCpIIXLnW8YDx0UM/hnWXYK2o+KyTrOe8cJ+BvmQBlVMQo+XbM4+lqAtUDlLZNeUOXeqgnujs
6S6UxVFaXTsu82O4Dcgs+2P1yIt0SAo/NGTdtRUk89Hl/CXwdxaVsuA2i4fsPxcujrF22zCU6/nZ
Ngpb4smEZ2QJSQUXQkW9/hjTv3kYv90Mxa5M7qRbx2yzcwjSFHJFeDONt1eBalzSh9TD6yCra6qt
meHXQwkLckZ8I95rROv7JeA7dCVGOQ08kQKtzk3CSAiW6atxL4UGkeO1HMZ60OspB95DMtHtqfzF
bdUY5mkzV3GkO6PM63quDql/czv24/7F8ntaFK99neaHUzIuIS+mmNpyYz4UWxs0y4v6r0YU+Y1i
Mzf0QainzETjn+hjQkVqT0PtKjCgV43HZmtgLnm+bz0y6YDbd5VMBOzvMIZLMe69f1wgRNUjEFbW
ZD7Eli7nAy0Q2KlB9Ds+EVRuC03F4JN3/aYp1v+KNGPRuEpgFK8G5A++pt2gvBs/2ywFhbCe+eCW
uFH14PIa3q7hNhrRvhHmm3zCvkOu2Y4H+sR4NObHMNMoHITPzZ9OGW5HNE9TLhFflvAPEc6NI+0t
+bcM9N1GWBrldFt2j1bBJPhKMoBFykXqF92H/1ZouSxJyeubk6BnbRQvjsqOgCqiDiMlQH/CIbZ9
iYq7RIfh0aOuRiUzLhqdnqytmN6QO+7fFbHIaV8HhfgVRckbW9o0C2VJ3wSyKHE8umVGm1Xci/SG
uo9GS9QvWCgLre9jhAg8h2u4YgV32zuCQaWfXjhAfsFBRGV2giieECZ5sKl7BDZCZI5lVCJUth9h
+XlYy9NRRnBhaIU38O5Z74XJxvn9930LLj0cnKOSNC/skRwGCet/Ym4oHl0F6puLZW65SBhlcoBh
wrfAa2t+TJN0aQ3SHZBzI4lTqQxJHbqbHBM6YaR5eF+MbPQzmpzCPPLhoEQbWobs5wKQ07erJXnG
BsIMM3kPP6s2rceaIT8eh2hjL4c+1ZRLGx37/xBNRlEB+Y45UQ3Tj/KvpyYBeDvnZ53rdG1f3+dK
Ulbw7qEtx1tK2F12/PSFfVHhaESHJ8kmj2BPdJvaQ2hTILJ3pfJM07LUYjpiNWEEtXcQ4ljq17L3
JPpAeVyBH46TK4RxDjLa3zvjpWPoAu6Nov74+jxgOjH54f35ZKfbCFcCrWAG+VkS/7BAjfZeYMUT
QvdrMcZsOWHf3uCmpsTpcfncPp7C3zZm07uayrL1pjrsxginRwNBKRJpbFZeRJ/sJA921AtgcC36
Og1bCAkFo5pUJnjXV5eyrLyRINbYzW2EoE5C3fWs0XsabPdXo5BnsCw1rD4zIxDpIIopMUpYDqBe
XPNUsnPpeTwb5vTnSuONGeaOGLMc1ukI33E+VDjMEXOgrNgYGRQI0V5TjkjvnOyx3gKgVdOzzeX0
OAA/EKGG0V4Gro4L/4o4OhQIjut2CjKatjJzM9EZa2RZlXm4baLTQ+0MegJomgOD4R2Yy3gmt4aC
sAdZXHqNNrvj2EjdGHFzwcH1d074tKuhPNvTQiZysQc876UfegjVXfW8q6rzzt6AuzBiBa8USzbh
Qv8jjS32Z3HWwPJxyCTy92UIRXOpXA5afVul+WZDV+u3qWQ3Yljs5B+OMqgMaiVkxRcL9gwgjHYu
kkpOPf+gPNs1AACNYx0agjL8r94A2MvhypFSwsAdLHyrowPztvs0ZGcGdI853Vsl+yiGlV5jx/gu
ZSwVg7aCZVfeRbd7kouUdrq7NqWVpcJ+LEmnlBOBxMWIf8+EfrHiwtMkBzBXcRpVOhByjJTdcWtq
1R9IPfZTX+xSlS40vz5e+XS4IrMfsse+KLSSiX3xNe3nYU2ZBTG+7OBVZ/aFpGUtDlc41/qKeUjY
beXCsgvxXB1rjGPkdbcV/igrrZ+HvRSHEluSZFp7rFtcn6WxArFcAjofcon/4RNdIx1MNcOg2Duh
/rMlhl/vGf4vLEh7ijRlzGW/qxkVy+AFz8i3u0c4nlsyvUVQy0Yw1w3NLTaH2BRQMwjtKLdn3BD3
ELs/nHfykVTYrPI9+Tf7WzhJjGdhgC0+4jOrUcucnrcSMdfbWQo0t0DyDU5pgWcHGreo4drTj+BU
wdldlMdiNn1CDqRPiu9vkxCHWuBvPNzxCjXxZqlcns+Zm+iucBwRhXtEVGWMWCutMp8vNpKivipn
3IjossSIqvM9w8VJTAL/wnlFGdNTvlQ6nbSNNDLMCXgvxMx9IFRmtQgTl9HXlT/wJlWpxr3MOoWV
v/vhrzn1bO72YYOBJmQJXFd7610aYT6C7oPIjruStGP28Xsknfisb6jO9rql/xgfzFgT/558cU3r
VJQUPqOd1VAUA/BLTmRxmFkF7/HOeN7itWYAMS3vKEZcdxjzbj4Tjf7/6/8vgix0+jBZ2Fbu8UFB
/lsO/5XY3VQKDnj5dxeAgHp3l6AUbC+TP+NYJt4mfZnSyZyUC8U9R68Jz/LSk/j8OB1vUliE9if7
ntL1xgBvmuy3S5dDv77P0ECFQ8poJ2n6wm62q17d140Xz4WFwMuA4CJW1ELnm/TIzgFdEaK2cqek
OYLXrdGtkTqsgeldNGygWBmMT5+f4AhQOKupCeyO5SzT+4F8ZtM/RYAxZXIBd78zokNVUCN7Hq7g
WU4HFq+dP7yBmI7ljVE0tdTCJY9IM3C8e3ADiGb25DtdLS44mx5+oYalvzg1CRUwbM9s+d9eNj7v
eNzEGKrYo3BsMtQuK7VZv8Kek7dln2gJCwSDhYX9msCj8hQ7IElYmSHT5i52UrVHOTtkAgVJSmc3
ZduUjzLaJdkT2pgbrS7DvDhNBgFMpvrAaf7NsxHZV5Nw/NRzuLPhWX54R9T6Eidl0gJNM4xiGR6n
KmcYIIjUUPnhhhYEOYr5aYTV787+hhgfSaiNK3Ia4SEWniPq9CSQgIgPFFAASliJpCyFZm0A39oE
z+25uV5q3uI02n+kZ6jDeDDLC4ZWCOE6FmcbYLllV7J0tQyr9TouZjiCU8DzF3E/jvc6HXtrdyjh
MH5P9xx6wuWOLOGR9JN+QbVnD7zyBW6tByXBySG5JfH2jYX15DmCB3AfCGc5+8LayzZ2hH5MI6ZH
ikrpGFxP2dUybxWpzqkOuE2Ci2mVbjIOT4bqnBsmN6Hgw/OtCOCG24zyDLKcD48+Xdjlb1rId9cF
ybKZHrcmCkS+IBDA1cOnrLtn580bCiYrLo4l4JeKkp+KRCJ/Ti/wbkScZ7HH8KpUFBehkWbq2oWK
zY9+V4YYPxLF6crHByMmTKfOmj/io850ZteFF9nhDyXzykBdi9y6ETUwF+3tyTPPceuUo3mVtQUi
OM4YCEgZTsGqz/jJ2y67FAVrZlpodmWoJ/rLxZeitYR05lGSNhiNituzJZOZPw1ODpGZZog1oF75
uhMmeQImamwj0ySiTRM8l3OAh/Ee9IgrbA2NEIiQ01LdAVZA9UANbUHOvFEvZsskQxgjDSdp+33p
ZjS9gIADV2NVeZNyu4XF/h4Bk1lTCBoqg7kLvrDuXaqRQtGyFc4DtDpT+LcdYXcsWwxK76eL/xKf
6u8BrFxjQezkPY87l/kxwsDrmtd9V7LQ5s/W+K5qsOdKfOdjz5iVK6X6PjnZmW2Sbz1m02sCM5la
i5BBRKql2qFJE3qkLkhtHq9bK+13F9sB+ESJw86tAEVUj9mKYEEUkiC9iNCTHnW1or3GlPmhS99n
5dKwUHpIc1BhQW5CbDxCUbSdDAlSztXDNTow3HMB345ZRnJm9HfakgBkMhPGO6Iel/RhDfeLAmP1
y7oSzt1xXwah3Os7G+2iWM2cltYxs3Pk/+Qq+MYyrvEpGT3OIrs2l37pGmKw6l714rDMEiRXIrsG
21FqR1y6qUggTLGmicdSPRgUNTM+uOn/bgjNi2WPBDNa+t17F46QY1CB9bGdAxJrfeLOzjJr+geo
xquL8MzzetY+7ED5qXN3STKrgdrnuvTyjNmcK8w/Q0H/A+57kbgopbo5nWclv/zjDMyUXgOEnwz7
IXnLyxQ8brOlmh8n2qY+gwG8ryArAzoaVYtqvlrkDoffYvDFQZvC0v8cjE+Li09GZmz/XZ//jGDr
+EZt1FsfaNkIKQXlA83IkTKJHCO62L+8Rq7JfXn7J+8gq+beCQ7pkaQI8owpcdfJUuyW5A9fSa9F
Vd25j2NEF+zO3vUJZeiemrjNzJvFTCbR+rfKoO39m32Oa/qDWaesuhaAFwodC9uJxJxmcIwSV4xj
wqiz2CNfudEVT5/j4cOEZe+7wxCwfougXBbRVmPsSLodkn9OdH1EWPhmSGY+nGjNnCYmdGIzBaPB
EEcKCVsCrCP/DTA2acdMW+X2dnUE+deHjAbmUQS2Hk/jvOTQX4Qts+XJI5NSQZiCm9d1suGl3Wab
lfhpjbl9sCJp3UrSylvU9h5WilNEpFy5Gqc+1aprAS+MjfRfCYHU0Glbkr1CZ1BpOJo8wqWPG/IH
fRWp0gHHMddOqrCA8hDASgPxh1LeH3uopprAoBUTZtQAIqX6DhLixPlFCJSOJ+wLssyXjSGUFo1q
cmsg5tlcuEr77K5eOLtXKAeJoA3KNJ3AlXVpg2bbKUoP+YFsDzSeOM/1De0DcnEAbcCnRn/W5B5S
NFNKANSK+j5JcdMBVu5jtRKjxL9TZ2uI8JJk00V9265U19Xb0XSh4fz5tVjqoFBiM9fe7dT1ju+k
1ppU8xiOJ2w18w/ehFTliBMsSeFpspF7Djw3SZ4HtHNs+zNJ0xIZdvTa7nsgM/jIheYebusjcpDX
s/TX5sG4H6ylyDNhhLILjOQSOMlC6Hnsqy0EU2wqrkwLCBoOlT/Id+SoANB238k/pQWDI8kl/Bhf
2MGoxmNLtM94FgNTozE4PiXCa74lex/fynQ5uz4egxJHFdo33tuYdJggS5R3DatUk//+p5Vv23TY
8kRB5yj8u1WcdXIMSSX5xPx9JZX7krs/Ru5E39ZtoEL2r9m7a6ra4GvjgV6wlXJRmP2Loq+Qt5s7
2vZsnH5WKJ1cfpnybcDtOMB8LVdQ2IbIryg34OtAwF5iiKI7qPDlxkBysF4piPIyJg6O6H/l2pN3
/QrjRS91mTei2y8XJkEBbLtEA/Bg2QcZqwaC/LuWB6mnbxNkC8m+BnFw7y/CyLoipyQcXC0dWhsu
nu+ysPgkz0AwD7aLAV2abG9NW5cDhho4B/0iVJt5cA+Tx2BX2Rv+CWX9uuOL+esscrdNEALZJLRy
/0FFFFNpAW5MY4qJDYVTTEtZoL1vdQktR5+1jJy4jGz8iKCHfvBW4+IHxsgy5TnylWrtNKo/LVwh
CdfR1jumkQKgynRMuxMmrRT165ebKW4GVI2IaWaahJwtMLR3RcnCf+xiIhJE4B7m39bzloGNfcBi
l8T8uHj6AFLBmJpZg4RV2xpf3H2l5J0hRyGInQ0EGcdnOyHjQXoj5Tvr2lPKHk+/twNPUJeR8fKV
eLxSG3EWD0PsEVIJzAKiFolAS4rCtQK8HivtA5lQyyeX77v1MLmQAYZp6tRYa4axqErhuGdHK08D
6tVOX700m/O1IjoMFZFgI4HbqAOST9L+5dzZU6ov8TOwr0OAkek9+UhInzbOUp+qUh+MzXRqmN4Z
8zBjXPpnKFphy4zH6GFGNz6kKQLbSL/tL5W6NK0JxcPdpDQh0CtbTHw/Zplw4i7F1uQluoOS0iA9
bSsNMc+Tcb+p/bkVqjSNyClOnnF8J7fEDnmpX97800apHUWs1WTmXEZCS3MbK0RBCeNnBpDagu6P
fh5+/NVNAT+a7R2j/caTDOAXhKrkVi1XQiSnITV7w/y/hkQ4rG5o2gGb1OSTytdwJYvA5xdkB4ki
zRHmIUeRQ+Fm9Qw/NKdMiE0ha1QuQyFALowCvhWDZSXsRnMuPiQyWlG5LtWw3GOusgwCdF6QfHIs
SOAWnBSG/A9Vh+PtuC2gcPfOHq40nPROs92lP5BxRZeMRir5j/fUOm6oH1Q2xk+4wg6w8M0IqEQO
GcSjit8ohI21k/+jdLLBhz/L706x/1CS/wIC1gcPEundmlvBX05VEBw0Aeb+Um45MUjG80JtWFDe
ZCb1jlmdQTm+8vxjPCAGrf68MVNGyyYcH0rbwX2YJSLlmbJ9oJkbSm81/9qsimytV8LJqrUE4ebA
vZGoHIpUf74Is5YGUbyAlq/wS0Bfj59uQAo6+b6HRclF7qeIMYEk+ETj1eE5qFG881eFZjnfcMPa
J9qf+/l8ONg7EOuOUqIgAE1NnvMQrZDpKzAIMT58d0hyhI34uOJYMLMSRfX0CjoSix5p5KS92oGT
rB1hQX33dcWj/nriVdlVKP7pIlYqRafwFZodbOzns77yPCK1nlHvjLOtFz/Eq3w3ok+L/8uhz2b5
I3+vv+QnF48A1kClJ+COAu7vwkckB2FZuraaLEGtk9HG4OgOskm29pnQZIrwERgjK2WQSoRwx56y
DOXLU4UMEeq8RutntFubRHbc4GD9y/Zkvx7Qtpi9a9Z+usVPCGYTUWkqWXeQMUWONUYvv75nSh3H
zGcX7xmnmqFZbGZrvi2sMtj+OzcHHiH9P7Abl9N6iMcjhyFSJ7UMKoUDhmTQehKyfBiKYpfa7aKQ
eUvS290nG0dF39O0/c5eu8YaYbkYDomnIxStJp/gJlSJtDbGJrVkZg4R/zdveyHYhkxN1b2DcXuh
1PeQHGw6Vdj2/Od1dcEshLGQlOI+Fvoe20R0++Mhh19tMlaB5DW3FIIbO3SxVkc0Llqdpf47Gpgh
0WRZtAA6Pd7yTN4MJWOEmvbJ3dVMGy2HyKJIukkkZRJMaEF0B2e9KzOdMHhKOiI/YdZwLOsAz8bV
v1Orh0QOLdz/MaZPhlvmu4tVi3oNC23AJrGOHo8UP953OX9FZLxtfJKtCNBRDDz5bxwDP47PhjTi
n8Y8Cc5U+PotlfdNs2Xkq8khRyGseKGM3es+u8SsRJvmMMB6ZK5vzK5ULt9vvVDgXyIK/B00CW6V
NFzitKA8MexsVPjad2htDum/e+fHqyGk+vYwg3AIbQulGLvx4iG3NWSA/cVWKZ4N+Wfj5ZF93Dul
yytuS3uLYMZzD2K2sN51hB8Vs3PZU3NKvrbXO0nd+FHKSO7RUgL68ppcanxARWYEU0cHHgLPK+t8
q2KLGqTHR/qRJnx0Ltk6zUGvP/YWMAq7SuJsYkwTu5ciLjLZ5vhx8qKAGEvdEh3UcYsmdpyPhevl
u40MgQ4s2fSt0YDWLYkRFm1A26UDZXgtWmCJABvR3Vc8uqZBNoDWoEGQlo3m3/Ri0pLjMGYtLoJO
ihJy3eeXogvzUkttPdE1PfFcGq/iobUrJtNWU0Etqn7xzaapPHQkbEDK92oznZIv7xFrccBxZLKi
l19Yq4RRPIuuHhlW5IEPeQE0B0R/n0y7+YbWzae1wR/CuUoYcQjauZmQ4NWnP30tvKmiScIM/UH/
mEdRSEHerzUnMKbVw9Gj//6+d5dSuaMfDd4K+EoX2ZxcEWPkelv0gHMFNQON91NA2uf7H1M8L7Ns
MaAFHYfoFyt43S2shwAyu70/6nvCORSmkfGaRzEf2ddpfW7m4+QxmZFYMZPX/la55apdVW8beg9p
TMP42jN9pcEzDKsBqJQo8b0Ydp72DljiT8sJdBjJGZTyFCkPdehgbOZk7OHzmKDflNH9r2t2GQn+
jK+L0rkjXxEA8mHzNk0I4sr7kLOJo1U9ic7D3Kr/8k2vdC3epYuYra9P4ejz8aY0ZF+7ysGYhXH1
lgaRtZtO+bnmjKwNwlkL5qsR7IuGx6YQPzE3ZyC1fjxHO8DNwXMvoktzWMe/IFzJwvwYdzoexucb
yqzEDTtFG5QkzDSXm18Ww4mLfvbG1GbvNcL6KFMrJEJJzYf04LtuUN1U4zjokYQJ6pCOz+MZJYlC
eINLachT5SdaUgDAohjDLuAjeW4QOa+i/lmvp/ZH7ujfN8rVU06iBPGfz2+FKoQgtRQs+ZinSO8T
YnRSqAyNoPD0fVJGMfp9mJYu/+DRMK72FYzXXtna6CharviMpqj8D2pPClcaG6bVEFDTEMS/Tmj/
5ER6Z3PxGHiVIQhFrxIoiLJ9pzFcnQnVzsl8X8m7xhoZZwBBQbD+ZttId3MsGGXFK9I4oVD+AqJT
mhVnPs7xUtbsDWimUT3b/AlDa5NrObk20IhRCT4az8oEXoh0fXjsGiExJf4MiivihhwIZI9RhHVR
wsjQeJonwsufusxJ4reYGpludoEfoZ/aoWhSvk/vW1tklhEPFWnqkQAgizKdFxSv2hTRqmWLBb3L
Sy1u5PcAgpOwyTBz4qclPHpGfm5q0fUwPY56Gs3YDMIpLbiODF9QryO8gKB+5RINVDnlya0VNfaO
/iDltzQ2QkkgtIXsiQlbD9lI3Y55/qY1GUTGPZP1mlRKCG5rNQAIxeOnRQWVvqVhEsE9sOgR7JHf
B8Ukoual8FD791KotqXNfTQltalpNF72WoqMkY0FNaTpI1dXp/mPf5C+WNYkslgQ9UVfzuYw/H71
6MxlzdEtmUr5OlBq2q2IYCXvFwC4by/4TlmBPV8+Wu8wGtNadRmoAPChuYPTEy2CyE+PaNd85nM2
XeXJ8AbV42GOgZxrs6hqGv+EzGVzdV5libU7oI5KQpFxf6Y3X5tRnb1pfZJNUJC6k70Lr2kjoXLo
gLUlVj8fwZPzlMHqGUBxqYDhjPpQ5GvkVknQIJTP6B8nfSPKQJXciOAYvI3wQ6BAZLHKwDYo0Tau
GBEQqVW7Nzg30OQSW03JnhZntpqcy0Kmu1SQkMzZzz/S1X8a9NiwPIKBQoZUcaFrGCsrSNgzowJn
7SlB+oXq28E2g0jJ5M5DVdpeUN6iU6ky7RvJoVUhZo36kYPrmG1pAGhb5K94drdxfHHBpI+57MlZ
MFPJVkjaENOL4Gt+1kOuz+a0/DtqmXERvueWJPIYEPYxQDlXMZw9OTxG6uhbCB7dYeT4a4rtN4Nm
faPYLxKxoAkx2y4uyg10bk8NiTbTYAvN+RAi+DikeAkyTgVC5snbIEEt/X/6/7t7fBa0G1j5lvKP
ZaXmsFNZrHY2b7jpnRReW9fWeNLiyP9KWuw/LhSAz02T9//paeR5dC17AKrwRVFLcafhbxTSQkln
0SWXnOY+DI3G8V38gcUP2Ubrz2Q8PYPG6WX3q+grUMJ0DpG44UUBP8J1UPSBJLP7fD2MOm48V84u
sEI2RJ4h5YAcxYYP2fog1vYM4ml4Y9CZklWQy8GA+QEKQ0kWLhcoMAdZCa+l3WLEdXJY2d7Q49Yp
S8B9qzmrJeC9RHjJ37qP1HIQveVvD16DbUaeNp09ULuHFn4fDQ6x09WLJhffqpfPodiDXhKEy8Ry
IvhNP43fFYIP1MgR2+2q9Ir6ZEt2oft9gXhjeCdu8PWE7OnKO5HMxdYkBD6NlKYmZA9zhkhKyxTa
RKPOQozMFIjaNsU58GMEtFljZANCX9ArspPDlhmGePiMceOyN1KrN1TnoH/L1vULDNkgKk8wKOMs
cdFMuGizwQ+RdTpG9RR+BKJDlkXxAXjGf0Nb0HO7Ee2eDQTxZ6cEkgXmlsRBLIHsD4Zl3qF0wfar
HvEBsfrIZndBXdduFanAK7iE2VhBbF6d9cNq6t75XxEBeLekIkOEAxoB6BrbnGBfMP0eu5cN2OlQ
wXjaIxfERTMkLxB/ioAogYfZxmkC7glJdv8iClwLBvmqA4jt/hGlsl0EmTJku8SKyMD1pBh3IsZW
yFQ1QDFt+cxGIl2uLBCCjMUThjTQap5KKkYaJ9TK8L3e2Bp0GKvZMjj357B25Er66QF8c4Af4nd0
tSfEcGNMupGmKg7LkHEg7ioaeGqsinvK9SdX5dewXKms6jgMZkHC0eWqwgwnqRqyTFmvIKz2TNix
/XqFQO7ZFAas1tPLB1pSbMI2QpPDss4eGAaDCj6dW9s54UqJyT92H95j5l9B8qY19+il1fAX3OwU
0IYoOnHUwQBRdE+Dg5jyIF8l1DB7ZWybgVAmnWfL81iRXxnLiVdq+biw+NZ/K88kGovNNb3IoqeB
B7HQozwMBQ9jM/uozUBke4jhlxEJjs6asFzzO38Be9CmR+/ojvYG6JGnGRZBht2s24MCdDEGgSTT
FUBkMlKdrrNTDVDYWzon1gDx3U/MteYLcH3f5TikBmVqKvb+fiDXRflbeizdi7GzEcJwpzLO93oK
SJHvkC7rb9h2PEJzlKPVanOS35N03X+7JtJD7V7+ItAlPQ9WY4UZO2bHcsaXPBrEQmCt71xmNkaX
rNPZO2WOAVfGBqApbIsBVq0VVwuBVbisJ3J0wnOtau803k/IA14/qAqqvFT0zKAqMC/eJ4N0drli
G2v7vQVKwLTuqVYLPi1shqn3lW3dzow6u0f2lV9SoON43AX9Hhoj0LW+ErzGfRBz5IBJy4hCqGAv
O5WgyfqZ9ZEcLUDE4iELOt2pxGnlcBMf53DQzUG1sEL4fQoPFs1MFZ6r/jjvVshTYTDetku7Az0B
dBe0RbqcnC6nhDGvP1X73L6PFhQLMyA7NOJDJNrnBWaaK0rijywbfKVJ153bwdqIhZE59zeGMWj+
15g4l/gSe4YZwZmXzR0HN5VE3yO5R0KfExEqibSKpDv8exl/R8ObpY7yfa1aLs4rGFuBL6BIePk5
aC44/MNrpeo68ZIpPtuv1OdwL59mjqmAgIR1AC0HtWQQVhxobw0UvxqLtQS31uaE+eSORpF5JgKB
YOPQUIOa81FMmCPqH+EE1g4gqH5zHeVpPuKeltmDrsZJ3YP5zKCP3T2NMYZ/RO8CuNaTfKpa5Ue1
MzWYtomgqEN3J4Qx6OeSIGwDerON35LTI6VVKNDyIVEsTekLElJJewS7/vXVXFGgQo3fIPuAq7YH
ubtBXWB1ubywWLEJ3ni5ESyxQbHYI8QuRAvcPK9EwN1iyc7vFaq1yOMxcAOS5lvceXFmtP8phdSC
95Aj2dCGdE/mc5Ffow+li/KZ8QUl2vkFC/ERxNp6YF/koH+WDtzUtxhXa2gfBlP7RwCGy4LOTXSv
inLJfycxriMj+Wh6ROgmIjxvaxF+X2EV3WZ9b193BQrTmFgucgA0+EZfu7qzvjGeJe1bPt4RM7s9
yhqZJaB01boDefvBpaAealZLDpQ+8hGZvibeOniePjXXkdNKTyAA+wEAsk5hRlHIXM4rXWJbAhF7
s7DOQVNUwYkim8Gp0Fj02GcwVPESBMY59heXBLJYP/Q/Ak1TLSI8ZQKcGYg/0bHb0Z4dU2vi8DwP
yD3SxisO8KTk2sA5szbsW6l+uJrd5okOkwavbr0i+GXGkCJ404McX4MNVMpuySguoOMP6ERgnWP7
Jk5E8296HF37T4rPGdIFDYNSGCqdeE5lw52u4h2pzMxQwh/xe3fggAP2Cha+1Ddae6EpHq3mzg9p
NPqiXiZWEuH1eGbuNMsGS/73EQahbxMOMcQHHxwq/AZovijfKK+CAcBU6g4m1JeilTCxKuUJ35hw
x6YbEYMGfN2WUU5F+BHqsTCTJ6nKCCteHX2yHUZTYQlZMMOgI+QzbviQw9QainHvkrB6nfuC0ZYs
6HTRRR/QbashxhtGkG/hEdpDdeQjnbCoJi/gIdayaojYko/RSJS1VqPaE3ZIYvM2boggyAHJ94s6
ypFNCevzv6xVydLMOI4DC2u90jF3EsPwJwMi08OHpZfHLU7OuAra1AHP3hLlEQZRxDa0120MNUOv
9+ETAbU04HZ61cmstijjsdoLb2i/aQamg/uvH/9lT4Xkk1L26o0h5wIRvbHODUx55sTKvYAkFr4j
wBCM37QxICSRerdpGpL9f5Nmszw6Rmp9C8EoXyrNafwOYUOCXUfn2wrhjYrxUQtyBKE/LIjBVXi6
Caa4ciJx603JNymEqveFT8ZKqRTZfuo7QKhln6rPWlGYEdUFbrGcujF+fHAjTBFzPrewXkELMXWq
/9JtWClvkTyPhZeVgla5Nsn9Nkg7bj0ycenkYH8dUTNYd9acs+Fnikft4B9pgdcUi5X2n4ZBVOoj
nnGJdVKLQJr/18HvkrbfOBEO/M8GofjPoKq5wjGsQs18sJ8D5ksV0G/iwVQDssORQDjagnhhm1yc
wWz6YPKnbtFnDkif99PIGfCxub1bXGJr5HJppLqjPuviAxfIghbTb01uh5wJtLgNvazBo0BQiIQ2
83a6HMkKfJFSyBgmZJ5KxJCGykDFYFFpUGrWaTGUIR/a9kR1zn80o++YzdGwSquujSe2uQCSWPDt
dbvHg+7ccOPHFFPmTTE1XYVa+le+5o2BPBfaDrdcVgUTQQlx2gaLCG2niab3W0CaT1I/a9cVKbMN
XkwUZuWNCysGAjLyVGscrLam9CGE90BSpwQ7vhpIulhJ3Y37x/1IdBzPTsYHKJumi9L0U2d0ovYk
obQEX2ivjSZt3uhql1ppXbLP5Ht9HtehGugKBCgg7/xmKbZpeF4Yw4bx1MQrfQvOTd3VvFZ3uuib
aHsAs2f5tvyebp6quCznOGcvFsZ3TQv8hW1DI0hYnHZrs26L4zTERVDh6khjQJGh1goe7UKZ+/97
6uallV80Cb3ujGq8+6ZpursvGodf+AaySvj3owSMW0bWPPra4NoRzwRPhr2GDVgA31xjYPVWeIKj
1Q3nDqD7D2SgHWT0ogdVUQfGZvUNr71p5pO7YUN65Z0M3/qLW+75161zV89hZlTIacwZOL6SkQ+X
ePsA4jezlUrRuH55VxrEd1CLLb1o5dqtULT46cVRE8sW+ACwJUvLZ4KoBMgpinZq4pH90UvJcrMp
P7fP1dvzYvc8OhIs43weFn6nAPJANfoeBIkCXeA7bW1SAhYnAAk8o8UhLVA4pP8h2pmb6pXsvFrH
Ej6uKAHXMxvuswLJRsUtAF5O2p058vdZgSAuokRE7G4V1FWUUOythq4GEeIUUAbsvfYhYGCt+5uM
SmSWoXfs/jQk2sr6YeWiA1c2ssz6UjykB2WvVpB9M+OFoOXvfQvmGpmnIrTudfxX0TBvT2sLe8z5
endpljb8faMW0tEv/vYPEqs2Aq0r23OGxWUrRjsMRavMrO4kYVg6afsSg0jSKRJGxTNO10tikLoZ
3LCZsNluEUONNpySUoc95n4fbbqPCpIJAxhxgpuQM2jLzDr68K8+ndCJ+s1ejNGQpJwyih+gZ6rS
dBmu6g/aFBYoikPZMysTeNmOBCI04tWxFfzXGdxzCk9DNL6tpjPcZFOnP38zXaNzJyubGSYIfZq7
IDQTlfm8231cj4xfBmCgCRJYf5+qHR5WrL2oZgxgII3yruSacSMLnBJP1yGWHaspZ+nn4ctf4kG6
IvxFkHxM3v1I8FaYzN+htKAfvpW4+e3pYhYKF0TEOX81Vj9s6mrsu+xF8ZjH5ciXTE07b2CdwkEk
LeDx6rbFeUuomLrMyjvVc4xZcUIUu6N02m0SrYVa49WRjpfEL3E87FnL9BjOSdd3RKYG6Hv+1Z85
31fRUZ92e2KlqVoYpa9H5aJ0NOIgNIFDgvq2m35YNIt9X8L2zUsm2lmU8d/ag54NSHO1+n5plHS6
G+u+CQfPpsWDOlLi6ePFZuIdfRsgShIIP0kgPqde97pSXGRwKsrGCdAoJnNNeS5DrQV/k7e12SYo
bcK3E/6y7EjAaDpRN9I0jt5BY8Gx+u1eFq+2Va5N0+z45FaW1JYJ32tl9unMQ7BRF39LleGA39xC
ARL8we9xDcoCFl0Ce7DC9iksFpr8lNaSv7TY+7M845z/FzUU/l6A2P19bMqUp92JZSogPkUMeh93
KRa5k4UTiMIO7B9LwAVos1uK7Zw4rJgC+Nn9EPDjGxNDw4/aZfUwsssCBEhyDr/HtAEzZc6lgBL5
fHJJg3N6Yvx/p4MrQRAgQ1s71zEPu+7ERjkk6PkCjiQ0xq//2nCSO+NUNsbMy63odi4n2PE2zqIj
Z2VkZ6dMwqAPx+7ETUQkT6CvTPjwC08X5rSGT7HHqHP+h/pnJ7jt7UdQotpqHatDkANxFONy3mna
q4zaGYZR833H8IXws7JBJkE1ApVtBTI21dRbIr0LVJXrGWxc0qzu88tpICKyibq2M/SXRUtqY3np
Q3Qy+JE91GtB+TL54mkBGigs2OvMxbagvOwHOpz9q1ydAvHMtyyramu5pdar+muhfAWxkvgJhXpq
3cV+yJihYZRhifx6XrdNDbo2HqO2bU+XVlunVmlhoNFE/G4ZmldQiDGy7XS5bsngl3/fMlpCewIO
ROdZ3QcqcrPZTy9/6ok4iNXy6qC3tr5obqNdbYUAPF9Nz63C8fPGgQOHaIUPMjIU0pQW0KbXIHQT
9ozFngY0CZkFhojtFUNt5LZ0Z3d45x8ptpDwhW5NkzkfgOOlBsYr1/xCYpIZPOTvsWr93/b5Zpp6
PWoW5F5M4Sw5Nxm3RmKXVK7WHLz2IT9fbpAiu+F0IQAl1QVtVq8kCaAEw1J0lDEhNBQTpuc2WWMn
jCTj+5hf895/fbxlPPoeQb7CfxrLY8CRegXx1cE46Nq581BTltikFQajXgyhY+4Y2MUWxG+HS6Ee
tzOGems3+IBSe4WEhaCraB/S0PK4hiqyhx3h7WgB1LP8A5ayDUm0K7xCcP+g7R3+hzvK755GB7YZ
qF9sU0a05yGlXUn+8Z6QpYpfCucJKsMLTCeKwEhK6T9fUEGtXx/ZPuN1380zmM62vSNdo6xpX5jl
tEpMhOLmuXB5l2rWeN06ztynU/zxfGO8NCuv036y41KB8LcgU9f+kFHRrc6wftvs9dv0ro4J0yYu
nSmP5uZFmA0TQeXWcjVN8jcITZUx0EssMORNnMr7S9o4//KMwAq5RbvE29yn3me2rA3HTLu1m81u
CkinhWHqUVw4NtEsofRe7DK62SM/mrAt1QoEGkTQaRtMybcA5gwobVo8Usp5D3VeM6b5ThWhmDGa
mGq0pCXeWZk4MoGTSGRc7jaEBJK2hZQNrkESAbsxY2tjCCqRrYKI53dJb9hB5b+IwZXxMI7hdT3o
4vV99B7Jbt7cVGMs6/Zz8NAuM+D9i7PX1lgR1xCyiXVBTm+e8ntX+ZylqUW7qKSwfftAy/7+8urC
netNYHdwNENYbuvLfd4zH18DopquSSIEOQWBL6ZaSgnzRMfwXCLwQvuk5Ayy+/X7HE5iskC0MypQ
uS3aa4Ptw5CuquxqLbgwN++FmkArW34wyyODw9PRwXY6FDsizIDUJUpATAl7aYITeiRUTNXYPg9q
VJm1OBBK21/r5GmjCZWUYAlaYHeDx8pphvwGvjRDtV291rQeQ4743MtztBTROHerdAXM72tWx9Gh
be2kcoqclxZy1ekpnTvOzYth4BXrNTQB6uKF7Eq/V82nwFFXLfe6HmrnPK3QCVht+KIJTfwMjWoL
u+dOIB7Qgl4wODdVhSakSk71/zUc4NAY75xKlN+no2GrAczlCmndkrak73w9C3HzgT8KCnZqwUs+
hca6+cib0mosMYxTvOrYjsm58ztdFh8XBbW/sNFmNpA1uGg/4WfkL85HOlvTsLlr+FawU1SfIwpK
MkC3pPUNDy88N2CYJO9XRDaP1Eu/qJwp3wi3UsdxtjkdxWU1JG/X1ugHWcGAdpJKW+YiGq5MwCRe
QJ9mKiRqXvJYFYQO26dJiAgg6OJXNscLWvLe9FF4schbatkebgG1iFMEVVxSTgLlb0Y001KQkNjb
DIFkCGkZGTvP94dtY0mwN+dA+i6xZQjkuurUepBdGtQTbZKl32m/x5eD2I1+pXpvx/wCNEYeC8kO
xmUbZtRSj5oZT7RIIRkafFyn3rLNrSoX0IsySV2136ZBJDyJJ+f3Pxjpu2EyUbbgVPt+gOhQIaV4
U6SMgM30u+lElnE26YlG4CSiJFOJwAP+QjPsXphU63Cc1yMYH4qWTGhFffgYdsVBgFPMOjeorIIX
d7upiG/G4oRRxsAo3bFN4zghwpwaVr/BjzJXc4FibXgS0r5jY3JIp5i6Bd0e7ZxnVj8eqLrKvMjc
Yb3sRGWxga8MvBa1lseY0uqmVoRKcAhT6KDYmcK3OyP1/xpjMXjDghZBNk4pGYhMXJgBt6B//c1A
VWUox2pozw6NCPYLYzGvB6vLzQhL5GsiJJZmnJR2U8X4O+hx5z3rHKaTm4VjCL0n0zIS/9NasZ3N
odjPYDPDDYEpw/apOa/2sxL8Ah453PvFCaKDMnCcEdYP2OWgktbkppOrbf2iggFXDicOcgB++6cx
oXFdd0KTwoKfnksWBXuZkWeaLU2dshwq2OSeLnHus2L8fEk4o4YVRgjQXbiBxGtkR3tgMzglOuuL
WE6KWa/pBiucrGV0Qrkwwat2dJB1J5WDN6vCJtcln+qwlsMDDHD/5Uu73uA2gyKjlc9ARxYRJC9b
gEmP2YNFzXOcByllgSiz8Y2RKIEvd+pZnx+5ybL/7JFDkZfAVuTxTuTsHwX00RDGmv6M+lsKMG1I
vXNgW6Z5PKYTTDfpMKrZ2JiyOjvVenoBb+T45Ojf56FkxFoSMQa1bQ5zQmYPzTo5Qkj0XGzgq9Y1
LzbZCRXrMcNmg5KkkoPPf1RJpgQAgZx2iqy/hUSbFtAHO7gEIBDgQFTMoI4CY+06hjguwe4TV+Ll
sxDLZ4i671YGzyHJmwS1sPitw3+ZyxJ6CEjrLmcWQwoyMUJlwUkBWLWFuF3Quz68qt57nJPRVYH5
piVDoILQV+ulpEUtMcdD7MHN6u9kwdrcEVe9Em5XyhA+TwGv+NKcOtyK4Z2LvJ03VLj1Az5bLsJr
PPX+p0fcelSNemH+QoHDsfnSlaWRO0rpixA1fWXYFSXjn2Uht7VyzN6S19938x8afcYXkihEFIhr
dMq0XfiQgj8a9/+gLTVfmXevlRwOeFcG2MbOMZ31F4Cdv5M1tFor1cM2LwCY7pa0+K6QHY0H97s5
owumbAdXbkhmDK7GlkGIyyD1/aG/x2W/zINk/mPzR007M8/kAi/PXxoWA/J7BZq1eVz4JjWwK/Xe
jxfK/7a6yA7LQujiputEAssR/H5O7IrlzVBJG6rbnUnOkcnTSW/PpO87OSlXzZsGvO/4fxoVrUcE
c85duwNAFtgqvaExv/w6Whzw5Pnu1hWViRm+iyYD+dMQCHJY4PlCqiPGqaUBxsp3UjHvr3lRHOfQ
9bSJKeqYGb8hpoaOQY6OSXgITKqyoR982RYFzuH8Y9LlGZltZ00T0dhZcB9foWc3aWQkuvGx6xvy
9/9ynqBUknvNsB0qpHlInTkSaSjWHBtsPT3ydZY7Kmd2TB9lNUaoPIN1E8ndQki392jIzBG8TOUF
ezemRuhWmuL8lin2td5TGJhVBNTSV+RE7qzf2dcHZNfUN1aYCvtmW97mPKIsO76+PPcAO/N0Zkr5
yIu9qnJwTeQuMb14Gue9mlmbHkb3YVeWCG8QMXnWPopSpWT3l95aytNSmAQnUppMR33CY43pMOHY
RfUvi+CRORDOO5lRpgWCyefrzF8wCWmbwDGZXK44Hgkgg6pHgELa4eRLuuGLA+b2RFj/fzLs9U+L
vp9e7u5HZWH0RGt2DKD+84dqrQ0w7Z5XA6gVuVVBoHPF6oBVNHOKgq+F+wSoKQIs+lBit++o+5lU
5etbagFN9pqTP8kM379x2ZmSpX9G3qifb9jLLed64mzU66cVoPezarXqiJlY7XNVzF/VuCaNC8KM
HS2Eecv9ej8gJdzfDKqxGAvuUdb9jng1Su9Viu7mmij44oEVLEub1hqVGy8qkkANH/mqT/5Q5RAK
Uu9Yl/NEPFK4d9OtHzZcXEOg9NDGqtEAQeWqxaCsxv5e6i4sEqec3oDWZrrEfMxAPY0rdmRpwuKL
grocdab55DawaclRZYLgtXZVgGcH6t/s3TP62VI6KxcOhSS145ZzqJx75g6QisPLlpbPyZ3cr47O
rr9hTtw6+/u0pxcxVoNQwOCyh7UwsO5akcu7fLrYAkMctB+q+Hj7DMdVntAU++/QVKaZ7q7ZcirP
HrKGsEEaPSy/4ZddNUR7cOOpazTZ38UoCb+OSjAZtjeqfBokxQDxTjs5FKvbxB7gcQuKsMqh8Ek/
JhWAVdw6Wrk+MNj9AEyrjjMVk8EQB5kPaW6ko+9+giSQFUqA/tZCLtfcXBwGW8NkSylX34U4AfdE
DQ+cirb6khHg577Ohxh0DkNK5UmKitseuOVyE6qWQPog1X6lYWYq1qjEcjhjvpP6+VjXiIn/RuBm
sr0hUin8y9u3DZ37dmhW0pbjVM50R03ACgUQJf583+AiVypXiz/YQzmFQMMSSMp34EYf3eayOHMk
ocXdQHMfsd/k9GMEQZiOd/HkmEahpUFGDp2kxbtwaiGI9B5L4SlS+ACdjDUkDTFSCcXU3NAQlfr3
QJjA17cqp3WFNGrXlV/ylQSqLLLMHKjAKm6Yiy+THV5L3GP2Kh5w5b28JZpYka43FOUB7gHiF59i
JmcIRWP7rQdMzZ8zpRTZ2f7R6eGwSJI7vX5ngO2euJ+cysmKZiiPhwJiGvqz0wzs9vvzCT83Aoae
c9R0GNZr9xXguM5OA9rjGzh5GDUpIx5nQS5rvQXXna9UYRpJ55CLQcxFThr6X/FoHaUmgQKcAWES
qUZ7eZBSiRf8Z7r+eNTMrzXQaI+X8zfgLfCmSQ6L3EjakcsZ2bYzQsumVjEAwx6/WumTCgI95Az7
FOnbLWaxUErKv+iM5wS0PbSmDHBJsyBsTffyhf4GNULcSKLIvKC//EU+jhL47Rh4e1ienf/Y0ftb
nPBEJVh6v0BDHc21esNM7/jz4KOYQu9Cigf/CdM32QV963cBXfYg8GJTq8z1+2ym/uDQbWl4PyeC
XWZN7DH3opjdEquvTdiYjfIXliyxujNLXD6chVEkT91Tsl+FtSmx3eGCl7xFo2t6NsVvAf2/blAD
Gn0X2lrrC05SlQsdbNURij4bGE/BHVVcOX+emNpPfKkC1BbspPqzHnUgec+R3z680BcsZ9zK/IKN
BmrwJ1DYaphFtSpsXw93jnkiFiUMHBwxe/TVFeuAMpbtRXWbvL518O1ZTGg+9yULGa7aqVqKcErS
3CQ2mUgilbMPTPdDnf9s9YTDpiWBSGsO2LANfh8MzKv+lqoru8WB+s1uQNj76lGT5HjZMqf/jpA9
GcmXJ7DpiBGCEErdo2Sy5Q8oZZL48UV66MO8N8yiNdxRHNA3Twt9VibZ0m3VmqxLJwnokyn2aj2N
i3Xj921Zu0SgC18D9kjI+2yXRPoMBLiqjqXrBS1f0talIbsj51f/q1wybmLbuYjWImKGdD5ouRSL
gkNOYRaZgrlOlLi0Ch6PPHyyShTbtj5k8pYuzYHQ5lP96pFuJ/9RMOJT0EfgoBQUBTfigj8dzyLh
djNB6IY4+w6nIJG8hwTqFYvmeyZNggg68nIzTiLmItVDbVIsD1StEudkvfOAp1rkKCHGj/FpE/XJ
Huw7cIMrbPmAx4cQ+qiHkX5TQbWwjZXcvZ7Cqd0IgyDu5uD4uFmDa9cMLgMAiuAdlLSNG/01sgRq
KFLma3X3UMtgEzwjM6N/say27Qa00fH0sv2ZYh6IpehK/WUDNINlpbjgVeApvpkYODgrp/1iiN8v
X6wni84FJv/Idrbw3gTxv8qvFmhrzHGrNd+UF2+k7tVFL4nR3gSmdjqeaCr9q8n5S2eCv2u0yLEs
KH9jMAlGIk3kRXdZQwGKA3OyBVOMvDmg3A/ega23JDWiP6HvZM7/KPWu4eDf0wrMp/vEleg6x7tI
PWAqf20vA9Z5nPVHp7xvn2qM5FdSXGUGuHjV+TeiZB+6M/l8PZ1xAgp8ccg+mQv0Dga2vee4Z4wi
Xfij7W7AprqrPkmCj3YSA2iSdTr2em/+4ujGpCAqaaF5suIIuL5ImSBNDy4qesPAJW37eZMCVICO
c7GwMxwIxmUMITFKsRCpwNd9EbZgng36x8nsZPQaCyTRYOr372FJDqz/6piPor9UhZXBkQc4VY5g
GfHwzF+GNaGefcNQHcLLk0xJpoGviOey4wkchS+vvACoTMwTEMyguKV5lcCSEZFcDVsLNAD22b/m
36ZmnpFq27TpFe/KL+0BYRLXvnw/2QGZm/ww3aneavVtc5IeQ16qDZEagZBIzOjcsnZ/p5dutx3Q
NH1Z25E+naT9VvWQPzr7+PursiKdWumfYBBzFKLO6vQz01fpOB9hwLMO/uC+w2KbvOofU82/JuLd
DLfIztGfRmdiHxc/ZWTLe9TIELToXJ6YeoXvfNe7XRXBeTYIg8YAxAM8/Bu1yWoNFhJJIX2ocr9G
3nEwMbG6GC5GMBgTZJ0n3S1F0ZedLaCT4+2VZ0Jv8uY8CIt9YIC3ESKj7SMkUbI7NNNmNfzWcZgY
OlFkzakvRqauVHwgQfJjBsyIkZk53ZLafupGN/gSgujYkD5EdRJwhDLqPMZv6CeWR+HSbyutNJdp
smtOhdSnNfu7KTjsK/NCkfNTKVQS/b9JZAkq89lgQ2ZAbj623t8iVAPqJCYRV9xbg8XIKfhQ2kbp
Arf62DVejLgK5PqQDoueqN73BXEQfYsTcEnI9/DaDZNVR/LbYfWXu79OdqzW74qhqVMqHjB+4wm1
6sqC9zEKEI3GuLBZtktvnxnU7ZzZ2qf0fzepxgn8AigFQHgaBlMl2Jf7uNXeOEoU3tLu4GFQWi93
lN3rzpUSxO58zwrWGOsNhiVF3E7QwPzz/g0qZr30ExXgscQv89+NIdCXp43O9r1r2sd7QjGFkcZG
g6o0HiUhiAgLWs4KZgGImJ4u6YynzvpRw3iMiokr+O1H87ylVr8Qf4HHo7UR7uhw6DPqAFUpHv4C
CjF/EmY79tZalnYPJ5vrhAcUFgwufgBtFJuX9vK8ynQ1BJhfHk/UfpWS9F0PsEdkhw5T6/FNcLj1
rUdyWiReKtGXNwGHpkh3oIIHMr74C75AFu5ztnt62G6Q8aMjoal6NSpuRkcxnC0+lCpBA+GccgHI
YnNaIGTl9PlIW1rikmW2kgQFO0off154ytuXPguerPm2JvwlmfZ5fDFq/bbcusq9j3dIYOYaxRMJ
S47+3/4mIW9MYjwTMEzGwCadzL/ns5NKcLVfdeS1Rl2BSsc7nbFZrez63/UsFimY02SqhdoiTzEZ
TVQ00v849TynJ0C27QLyIZeBa43a3bHdnUDgHd1MsECKFgt18FTevBvUaQ2lTP3ClUNKq+8SL1nO
/wtGcsaibXbam858zfdpFzSIs3cyAA59cf8kFUXNqZ6zht4ptqq7XlfBUPYqMtAt9C25xvKu8+In
XHqegKEtCx74pkZoeDuxVZqLBCk2SBJjNeThYOwYUvNW4n2I3WlCkHghyqH5J4D2WFZtkAmXMp3g
dJLCqtrUy2SJlnFr+B3YJj+dF8a8L7IRut9m7zbJcjv3teiMyj9HiaP1v5broEjMHtuNELGEAapB
ljZrdFnzrIJuNBwrrOlZL8ioS0Hxoikyn/bnyqCD8hLcU+DLWmDpSYG0PyW+vloxq6ztr0xsZKvP
HJ6VhV8rHjwvIam+wim5eaWxsxVzXjukXWyHSQTDb7t59KKM6Eg15jaUwIqEq4KEuffTwHMHMXAh
+o0ESHomIkk+DKzfSsz7TGHKqhbsUWvkEiVlMwEOAJx0EDrjcPIeHxAJT4d2crODu2t9DBw2ymae
kibTPMhKUJ+A5rR5PmAhqibzlNVT9v0iUbnmd5WGBanztEBI/gzB3aGF/6xJR16Kh2TYHySSwdAA
ogQuDJpKp8QY8AFKA5m/GhilKgYfLhmxsox+w2HKPz24dIWGtHnKlo0HoiSJrr/yKXk/OjJBEhvO
1xSj/OLe7T8Sr60q7PN+wXlwAxCyMmGtSmGe0XeUdgoaPUeotHSV/IKIrIn7CxnN2XYr+eyuZCYp
LQW+nnyf4wrEaUQdHS7iF1OvLbvblUcsztQ6bVzTh422txovEPlYYlqrbEZqOi2QYAisYRVJDmmc
Mw0MX3KxJc5Wp/8RU3lx+v+Y5Avinn0Dx8dXyy8yGuYU45ZA+yP+UoNmhueeNtgi50mjzVSlXqG2
GNghahBBVOnGQCEWZfPXblRKNlLAiZ3+4ltPCmq3XvQewQoz1vdbC4rxt08vEE7KlA6gZ0eKb2i5
0tyHjXuYFcvcmeAquOsyJx9hixlwFIDJJYL0QXXkkEKUldT5+0TldowgEcxSfNEErdO8K5l4K/Pl
eNbmPnh0PWL6EsmtoU7B7Wv6SDCKM3nKsP2HU5j98VTwrTcvkOhVuBG8sRWGWCnpfgz/Agw0+/eD
iaYXO60icspfr7ROGZmtMqgNn9A2iMTCaSz/zUwQs5sWJVK4yzaamR6jItIHf1x0IREK5K31wcvr
L34dmYqA6KaFX4LsGfUa2pT8OKoQosGGKx7Av4t5vrtmPfFUQ0AR24KSviQoYwjGGOdz0viN/sW7
bhqQFte66JcF/lQlRXNDJmeP8cs5xYvcDTu7LrdJrJxqF5u9bbfH+MLByhaROjkQOStbHDub265B
lFYZsSCL+NGRh/TcPSDS8xvo2W1fpJz0vTDGm/KmZvlo+cUroKs7fY1/djhyUZAMvGrj162ZLPQH
0WaAus29cNpQ42fXBMxesVLGP9/y2FP3w9BaZnRF2YCpr6TUG/jhflheyLcoXkpD3xLfhzzTI7xB
sEQfJw/fBq87/ti+tqh6raoMbElZ4/RKwR8dnF3HT9vlkcS25Zof2ZyDLgA8316LA8bnAWG8uh71
NbuKlDoHJj52Z2bqiu0LcB+qLMe0sGFpKL70Jwa9Zgz6f9Gmn9Mc9co3EPua6c4Jjddc9UqVaOQt
7TvbbCWehFI6CxpaSHav1itlMlLfpBf9CIx/A6VPDV7lQIbAqC25L8mYnZ8nbKamdMIM5KvCqA7u
dFQHCuFGaHDs+JnoLNWN/CzczY0w/hX/TlT6fBKaWEb8Y01tGlT5tzCPhdieOCGHYXr6AOstLuWC
26s0cs1ZAKL29v5Vdw33Du7odwJ6PLDiV754pjslySW7C2pWzZYRaeHpxv+LyMFGp5If7fGbU4S+
p9rb8WaNMKELbnX45IJWTB2vrqVZqpM0663bIXD0EPtBLisIGLdGZ7kvVx6rNZchX+DyeWNMERkn
0ulY20dpXWGRLXU6OO0CJ8od+XdtZtSEGv26ENi+IUEPCOpXrnrcjcaT6cfa1wAJisyrGS5TC+U7
mYxvbyd5xu+H9HKNrF/lvXFM27Oa6YB1eYkHw0mmJSDgAkUjQU8mjxCufJEJYoqy6cj/TUwBUfBu
0uRreO8LjHlGX3otQwfUju6YLuAinekhUo2d9jMSv2JhcrMGlalldQi54AYa3fNPAFmh/EeDjS8n
IF9vR4ncAvRomG2yqv3A/3TM5P+EHtk0yokzBu+j50yQCX7+nnd7OTyogAB9gzeQ1mrwko/lzXJS
w5wLMO+aLp8kFAgX92taDFH73/BP0IL6MTGwxdGQCAobH6Cq8Xlj0tea/VvZu3umAQjDDuzIq8SG
40TlGfHT5aeZajzSsgqVhuF5bxPG41nQU2us3+YDKnDLhU4c7pCEsbJDAlaDEYX0a8UWmdt9R9BF
bZYyNULI/T+da56TB7O1ghwPjjrSU4sl3BA0Z7QFjpTCKgwao8RWC0YMYzSUOkzUcOwGYDXnvPDv
7Q4j1Jy/dtFeOSwAwctkTVlGf4RyGqopt+BqWLf8NP56X+blR+M7NFjoYEvWJ8wGeRTHJXujkVai
/ul/2HiVDys0IZRL9H8Tvu07YJdrWWifhb2clr/8LUB//VbfUzWsAZnRlI+OaY11/MLXQkX/j3ZR
VfPVIJzMc8kLefMStEKtBSTAnTCDRR1d5NzQGpcwO8S4bWYcIL87UJmEBAnAdFdG/GIr6JBka2iQ
sA4TyxipuqZcxu24rSjSP9b8pYRfdzE9eCcp9x2hAypYMPaYz+k8XDvC8GPGQzMOubCURoRiiGCt
x4Johz9wW15Suqsx99/ZhUpTpSzOKoQR6aS1bL5ffBZmdolRUVQInAT9Fyg1w+yg2HteAAROcDnH
p2/9OhOFTW/01CLJhFbHSqPpmwL6KRxe9S9HhLDp0IOczQGzlwOlGeOx1ONlPgaKRNY6sKOUJJPI
BrCB/lTcdEsjLbQLPGcmLKQbWyTzBAz1RilBKTrrP9U9qWgBOBKwcpx9c98000JWTAvEy4UemrKm
a17pCFN2mFITN5UjhDkNtBulHwWZN82hXC+9EV9FadNdl/7TK6y6e0Me9+42+iHNfXgx+FtdjxQu
tYtrAhdrmZCNUkcvBzzgISKr1Djdti7sP0vQmAP7mXEKdcrkLeOTvmjt1/y0F50sa2uKGa50w0OP
QzqLxnCa7Y3GoqLtNp7BEozYSdXbDS1gDzGJQZuZWMevO6Pym8She0MLtl00uPTzjNspdpWmBy8w
9nID7yyYGSFSf/ttDBymrU18CW6c2nZRPf2zUbYDRScGibnEilg8tTLPRedIs9GXf9/mQkHJIzWL
+WEUzd3r9kta5+LXnuiJt6XbhtxIE4fpjsAyBXCYeCmGURQ7nHvRF2RkzqeoODAKabRmhSF8TK+D
Wx8DT4j0j/vK+/H7C2QQ6Liuor7d/IgqQZjwRIPm1MYEuf6qpSKd39I8ZwRPxcAROPDzCqeOaE8c
xRmLq5k0K0fo/6Qoihd7dXaY9EGFYZOIRdPhvpr5nLwb3fiE490jchLAPK5zXy5OZnKU2jWWjys9
J5SEozfxi2NgUj9iytakN4NaJItjyOzYwODZImOlnNTaGzziGAGmDNYY1euGjQ1nsV48klV8rKoC
T3inSYTTOko6FurW7ge8VNZKPXz+FZsrI2ZKmUjwL9cAtcHwpH6DYrXW07rO1nro7fP1CTp6b/rT
A/leT8dAk8QWDXT7gCtjMYMH7f5bU88Q0mCY2Xg+j16UpNShAGCvqalZOHFFfQJ1R5N5Oe2iM5Jj
FhghjOX1rZXr3pD8yxEvgv61Jgu9h8FmFk/X1FFOUHb8Y/Qh0Kd6HselE50WL+V3rIzQBxt8sZSZ
Zare/YMB+bTS8iq57nyLg2jJ9h13mhCROBPspkealrB8NBAwwi0J2W3QTnAuryTmtMqbA0UOIBgt
FNjZD23/7PHQGyDbB8c2pifNypgOy0RZRn5KVcC+oceawd4HaENVb/omradUs28XpGySSbs3HahN
ykwmWnOnS7QeklNEalM+r+UPqklxzUE0hdU5Sei8DdKo3CmVcvWRC/F2/MJkdNtDLPo+npTpGA24
cjToVm3JBG19pColwaVObhuQvj4UpssBRz5wOG8MbeovxhyNKjejaQwEfm7AOWZMWDuFjxnKQryO
o9ZC70lWPk+vPBRLYoj4DJzsgy3ym9IFUGoWL7hogU6rLpMiEpg8cDGxKpz7ut1cGZI8cLyxF5dv
/SO0GIsqdEOmF0ZXxspE691x4rEOn+WtXZHGHcbOfcSid5CgREZa936I35nuwB8KwOw7Ufy/ToMv
ba4ciz3aPluuEO+k9Rsp7p8ZzFJKKp0g+DdUWUPfKp9rXTz5ah0d8auiziiYCj5ICvglKmMXFxsL
ZAsuihft8Qq39lCZJjLCCbkQYRUrWRnC4ISlvSKPPiHizq7Gcju11Ar1PdYwC+rjrSUBCuGfqt5Z
3B7iG0E5UgkCTWzWJgi0drAdPm4qzR+/e04HrKQIQZ2Ch0YagHZ7dTyipgGW7yLAmL1vvsJtwJbf
9iEGniIhCNjLY02AoXG/Ygq4bSmD3uIybg88bjc4qT0OqxAb+ucH89gG/GEhm8xgTts6DQt/tNij
mWqGwHD81xrzbt6wnWQnwJ251EsYQBjGKEz7QYtr6+GTQc9BCQO+oZSadRhxgbx7MeKG8GRHAPq/
FFBBzBrrORvE9BQGbkurAhs0nY6VzWpHyNStBsPCfBI2vD+pTS0h9ymru1yG1ZDm+dw8oemVNFo4
wXnNdWs9XY+T2SAl1PXq5rE3BEsQYT2BSlqMrHBxh1Y9j5N0MmwmzI2uH4lNzQ+JvTCmkQLdZN3f
vuejm1kI+oeZdZDrKMMFHWgb0KXSMrKMt1gz2j2Z9mGPeUxbfrSb01837IYy2mRZehXEGFs8XDoc
qVMgntHL7ZTDvvpI2QdAi8e4eQwsCgChcm0TaVuYoqU/lpUocjWhEIsbkRgfmZ6BE+zY65vWvyLK
l6ytlAxvGFtfxfy1m8Ce/PwuugQZFS9KMmx3VZDX2tNp7IHOIgy5v/Bz/48uP9WFKypMobJAuEcj
Kf4+ctbNsBo3Q21AxHnE43mWUb5PIh4CIkc1jvC8wpoa8ROV1OpVswU5CyXYW47/N4yDeBQ5plNu
V7aWWZFbWw/7zGWI8Yq3w2YFwWEHnr11sEeDOH9jS/7oV76GEay6017ZMun9hnpX9iRaG0Djc5uR
Ggw1VxFTWxwQT70Olnxw0jKHjVEasYkLKzkYw+IvDB2r6bWYJqhfrBhel2d7j7Ir/j3qWT2qkGVZ
S2GEa2QNGqAKvUoty4Axc2ksoyB4zv/xnnSW3eEkzCODOMpv5ToyP9ezBYB/obBct3Zopt/Osm63
gsCoVLWTik+g7rrWxGMrC3BFAlBm77P1NECGxYt+eAySlGoQ3Z9Xpd0DTLNSN9gmwhx+3fTQ/mfq
A5vmKWDEkBOw9KSi3B9rk1jW0sH6R5zLQvMwczDEpxIImHjmSfb5kaozwzHNUgPZAvzdCcNLBZLr
WKymYwd6OboP6+P8ZK0mUKIdbzcX8ez3GxhFriNCjebpp4pROcFjlr0vmWtGlI8dOSOQyGlkr4tI
A9xMwfky1ZRgtfLFFSL6alCfSAfoJvBcF0/JTD7d8ug751HZx/LpNVuToXLjg8tM/todKv7q2b/h
YPoHT0lLR8uB2iuXJds6FKctnLNdWUHZqZBwApBRoz/LeXD31vPIGPfvbG8E/5HOocX6+WfLk5dT
hriNUFCOD89yc3noi28FBfkpFARsBgZset4alDoj7kmthDLq5yMVi+CID+z7nfnQcMSeuxKx+lRa
Il+0ErNpWH13kLM0hFdlEomIrWwWwLAcmucaroPq+KW5rApYsniwAvErHqav9kS7EsjCkQ82T2S2
N+49eNN200Si9mHo6gvdtFFcJPBDhGdAE2zX0kDMSyDyKVXl+7axq8G0Cf/l8e8HeO22ydxWeGfa
XAiVjDJdPDypbKprOqZaKWAhC4l99IZreRFDrAmezvgq1XqmBejpdfhy8oeRTCCGG0vVbqErfjkU
H7KNz4qrD97If04c89U8A3lR33HF6pT7V5AWtSJMIztFH7UinzMRRqLpWCSGrKxtC0tA2x9v7kmt
ioramCGHcU5XwC8otRek2lTrXSBe5586939L9aa3B45lIOTdhqhQFBTNL/2nufrg3c1kG3CdD99Y
myKe/jIoOcEIDFHB9vqsvAP/9HEPKJaa/Y6JA/v/Xw7TkYxTs8VmmkozghhTaXlBrxJNdtS0nMYS
1Z9CLEuYaCSKiJQVlmKFsXo16gRq07iRjoPGh+rTUzFHXCpSxEigRMgwvkJf3J4JV+Rcwp2LTB2B
y60TB8DTvxCZdujDqVoDtJN0AI312xVAhtCUdRYdjBM2HIMBw6mmi2amb46Nzq60jToi6697nopz
kgPYJJE/7IX9ChbHT+Mj6Ec2TOP5x4nbo2SERQoYkgAqDhUCA7QkkMhLFINnr6WFdnikOrQ+q0m5
Ljwsq8lbsTt/iCx25bpUpK542+73lOLqcGknLVBbKkz9cdZlg0UQAa3Cs4l1btkGowvDc8Sx8Bnt
Mkmc1KvjlGwsqrDwU0f9mCEZG6Md7B7srnyUOwRGNSoCWXS91dFMMluKuMQMScvD6ZyXT46foIU6
5rWfVTFH8aIrFi13NPfoUubNrGbRfWf6ZnELMXupqUREKs3h7FRVDobE6pX3Cc6rGxa2AfnpHWIK
DlPZX0teffubITCCPRz4bGeWRIGyoqHL0UjYuL/XaUCH4yt0/gjpDeoVsNDg46+iNS8m5YfjH5WV
ZIigQU7Q3eyClil7vMvuYe7NyHZUibvQqzn+cZ194MeXkweTWbEgy6NTIZrKMt4KATO0ww54cqEP
LzOfiCATmYBRR40TNpNrT6oo5NacaunWf9uknE4WhZeyQQNPYCs5EoZxt/UBjVYPCFGlOSLyR8L0
UoAKa1tAn5CNY36bQ1jAXWyBT4fidCWgrjGSTn0IJhl8MwvW8OBgY9sjGqkXwQExBEwMsK4WfDOE
DoPboGnvsvqBkr9mMlmYsex5kW79xdr4IXQQ+ql20lipNWDS0232nz+Ln7BiEQOYtHlk6gzJUVbC
QS2sKboHHP9BO1Be5n7GkFS05GuVLNtNMlSfsItl6MFXeDuv4F5YGwzMxgfJVFekialHVVqzLRuY
ZIk2jUHN2ozeyt3KX4o5MUfkXfF4fgv+ayDhthrJP4kf/G61Z0aq6T/ubSU/TDTlczLHdl1cblkU
jjZ1BodCS9onzVOW3FzWypMRfUGGH2Tyd5/qhALo2t1s3HSQLU5lpwlDI3N0M71JQ1x5yclnlwtU
xfmPAeRnRK307C1vqn4UXEQ47w4C+fqwOYA9b0CPLn8kaCKyk5HYWYYwwh0P1HnM2UFrnQkox7Yr
TaNj8Bkc4ZuBCS8JWrTX5odB6sle+/vZmnHt/CEBGG8KyZ1Q5/h1aykbeggOscjGomN2+OKW06ME
nDWB2GeYuj41/R+g31adgdeUk0mdILGBHJAYUM9EBy7e9RK+OE12WCOHhVl4rCgFJbBbCXeO3kMl
ws8uaqsHpf6nqNHmSZZXm5CSarAf7IuSO1c9r9MUNxtCnCzVUb7lvvTqLmASrb5/Av0GBsCfCZpq
XrC0PvG3cnl8SJoajfxhptyp5d+yN+MVaO8JGp5X3nHoLYWulRpMP2ZXWEeUFXtpst6n1cD3OJ/F
2flFGQnHsCpQitaWNRpZrLYZX8nuCtKC8PMhf35fEq1bI6cOw7srwClieqb+XKfutwRbGBts7Lb1
K3vPwp0oNXSLUuHpIEAEGpgiiYNnGH42EJnwFXxJmFTqagc83ZXgpcZSaWWIPPBzzXbB5dJnGg4k
I1aTqU2wzwaBskwQsFw8NNW2mT91Ls3Aw4qnbzGli05nFIVqHKf6FdcbEVirJrQq2515+F4sDM6B
7C+oUBAynNTavoUbdfpMVsflmAv8H/G+nyRZ9OSFVpCo63RpVL4QNcojW0q2sGUB8PhHRA6XHNCR
JfcuLAuIYjaM3RGfD3xW50yysdrbzf6NQfB3/I2dpMfKgo9XeKuNMLGdk71U43xhneYF39dak0Xk
20tcQz6kUZtgjRxgGkW+39RKR5Lh9yoBCV52S3ow0tX/0+BP8WE2sWhD/Pqikk6+l3ti3CEXT8tm
xZA/9wxGO3iHgogfya7Fg/LBA6yh5BfS4QR5XbZH4jzdvouiivqbFEn9pvTl5GC6vXftrshxlOLH
mxHO0YOXpPXrQKxDyki/M5nmiN0G87fODaDEttWO7GSsy2I8q8bZK34gpabrYaMHij4srLYhx26K
ljdSyko5peAluXUgVKVLbjR+EWvC1QiPGxZJgZR4h2j29VfcnAJiX0VnYDb943aa10ccVdiDnrYy
mCBx32nLKXdAD8zkFCn4gcpFVDlUnNpfJMn4TN+pO88BnJ6MIxttO4DXP2CHA6BPEHH2V2VH3pjX
1m1j+QMlRlZd9EuOngjNUPy2Rqeqtgzq8GYfxwrWTrKHefpbByGkUCMxO9HLR/chbWYGfEpz6aoA
oLKjBfISRQ7TpsEVafRX8MTyLa3SqS7RfYcUMPBgjBT4pvC3SEMMbXmFLbWCfXlp958sVdKlCZmM
STvv0fCkOUbw9p0BTP/dbh1e2T1ZL7Rp5h5KoE9yzcOtHnACx0S/pEHJKcuhLD5gKsGip4L0WADJ
QZKU44m8L/+4GoZLwOHHMX7gkhZ/FJcE8gDKvlIrgd7t3wmUtn6gzLHKoFDb+wp5vug1BK0TKUnE
v1yVjgqyrHSBmsU4DMephYkhuqKR9dnY1DnRLF1WgM0gZNbUnfDfQRzQr9xNkkCY91sm6we2KbBn
0Xh3JzJ3yJ+raJcU5UXnebPhZa/98JDu36WIWzNXPqe7j4yFV2D1IsPZcagXQC2hAUTmNzquBsFQ
4+JN4ZAELNBsGcg9iEzsJLlFHTmILz/HG9EJ5apyakKAyPVeHg48CA3SKHRvTn5Yi74fXNl9aHuv
IYQT9FPH8qYa+NrvACbJaiBSaWlCWht/2goOPJV9Gy2YC06GS88P8eygoxG9niRViJhI6iSCU3+5
sxNrtJfROf2B6EnYaOwh87tXVoqv0NUv78i0cFJ3zPB8N3NiW9VsQaqr/xJG3V6MWgMRmwYe09Te
F9Aw8QHBdbCd8II5SByES+IzQVNIE6EBpj5rC4wra4tez3Y15JZUnGf4b4pJpREoOjdrJYsby4db
uLxa2CTd11psU59COPk0OV91VqHeWzWgKZjfuXSJyPTUPURmQHRjuGQhdUfU98Cq54KY1JJO8u43
igczZ3KgG0ID2OfigxJ7WIGl3z1LKLVDXEgUqNmeSMYwTNMvleHl7S6sYdnX3aPapfh6W3pjAx2Y
ku3rPp8QBk/yujD4e3H4N5MMBTvbNwtrRSlw6dhOgFxZbZRJNR/fyJtjoFPDgfdRq1DZyMvSUM7N
ccGTmUxyiekeACgCEZqqIbk4qEGy6P0N+nE+1cZRHjklIfyG5sRoddqaRW5vvs8njsuKINtphcLS
8aPjUv2Ii9LKuDmGElz4smUkSMwDzp1CXnZYnZ3359Gfmw/2IBV118ypq0LSwR3M+25lCLdZiXtp
YF72s0rf+6R9q3LDHaX3vrtkTal+vsF7PwMeLlZ8DQB62XvmnQIZ7gcRg2ZVQxHaXbcT2pHVSlDg
iHBYdjkEfG+QhdSg7YBjRQcJWkTlPf4X9ghDAeb6agNBSdTkwBAYw93CzQZoVxAeBI+qQ6Fl13LG
sJ2Key6gMpL6jgecXm8mGbK7RKSxsPmguA7Bevx8bq8uiSVU89EHqFDbGjEgmik5vTv8W07K4sJB
tKaOT8Ktror/ezRkdds1XQ4fLZhaULMIIh0H4CQ0QOj4+iInG48gNo7aq2baYHvDnhbRRUT4vkRc
2VLiTiCu2QspQUs3+ChhgYcZAjZBgG2nI+eFrSDyWOMFYwDmIpTDg+QpFS73mjQeftmaRfXBqOuM
nfDHohX8GmW4B00K168haEA6A2JqIT9gt8jMaQKON1DTdaGeMHuJMUexd7f6KGzWGnt3mPwfLARA
11XLkrpXofAMc9NYBmfkqcIE/9DQQGHqm6NglQJJksR0CXFcvdDF+ydBjmJpieJoTGJXU9/T4mqq
LzoOMDnBHuPw15BBUyb6pcQ09tziZaLzPwEm+YxTXtPmZie/yz4nTN35gof4L0vn9ffW4O4vHgRH
2lYWG5Nev17DdBsKV/OyDHHQe1QKp9mjJC+SwvhdVrtylzINK0FQhF3j/aSiBvbSff3qRQgC3Bmq
HjrLdnlnzv6dRr5mWEPDcfL/c2x7MP/69SUKsDLFPL8NGQgPYdEps1OhB7KwnkmtEpCI1O2zWxDC
yqJm/8wdQhRRTmV3apxaq9U4BjkJH/qSUL6CpGFLH3BxD6k8aaguRlaqANI8/AOBUjJa4+MKfru4
QoeK7auj12u7LMociuPVbGzZbFyh1gafW4Rh9AN6LIjajWOGtVqTi8HBLO+gqHNxlk9kohAnNs50
+JPWBuYkBiLvmWEsxPNbXTKLbBQ94ck/2utgpzaXM1sP4Cy12Wsuc6znWtStVadnMjysvnlNWjIP
x+nPC6pInnGS9x+EFRKKjE7QLrfaJiwkmQbBjisxvDZH83lsenNUZ1IuOJ8+oz2AiWsVGl9nRaBs
GsJkeceCyG7YFVBpDt2Q52PqafMQtscv+gDRaALej5fN9a+Rz1oCK7IgySANJ995kiRbrUiW4V0/
8jHP5/lX5zutnaM+Q5AgWYbr9WAl1AwKa63smA3+lREj1gQML9jHgIZxoM7biW+a32YX4XYwHzHB
Tn7wMxeel7DdPuyRyiCehPir9RprkvtAVkbZAe2KUHqZUzQXJm2h8OZW+C/z/jqnZFAuDMbwqry+
aMpXM152NeaBNia17/I4QPul+Km8qsH/nPc5tceZ9mj9BSI6GGJKUxza8VjfBsa2Bv1QnWTMq2gN
LDjAz4utvpnh9g95MJq3yO02TCV9R7jc8KcoHkiTCc32w/mLS1H6KprC0qkBWHXHyks/i/A/vDta
LA0FbpxhKiPqRcRPTKnLqcNZHccUoKQwHzktP+tdsOT9rTElHMRQnrY8v0jQtjCFH/veeYtfl3zH
VDJXahLWLc6jFyOlBDqQrCQ/zr5W1SUxIjlkJKQAo9zpnnccVEzH+SsAHk5WO8wlFJ8XvG96R0cb
54wJHyqvbfQ8y9PzBMiDmAnttvoW4tgHl4s4JARV/c7929iAn5tGz9T+SsmYFYdzQlh+SF81yQoX
KP+StTh0BPspXyE+Mqu6yOqiOCgfW1ika1lI64+Mohyy6Nr60sJbUes7kkrvflTVgLx8rUpDsZ15
FawXu0nxJh5QCMs6RtkhOSr3sMgNk5nYAmpTDSN2Z6h8Nzx3gRQyip20BE0Uwc/F5/z1oq1r0+F5
Tb/JKFxIfLW7I4rYZ6cR++4alACutaQi2Ek+YuTrpEgghmACSnu7NFF3IGbbluAL6d5Jnmt9cPzx
Hic3oDYrlqDly8FjstPg1RxJwJUuM5nN1zU2YRz6ds9V8BATgmHkWEyEp6VzK7vRKzqChOY6i5gK
Ay9UNf9sDYax4EosdwrJjFNUqMJKTWYYWdoI3MH/MhgJatFzRE1SlmdORy0bdhEcMxFD8JmhSuTF
cYXpa5/bNANzxMp4xN40fnSbkOiNgeT+w66OM2YZxeMr5Jrg3RxXur6pZEqCTCrvJHml8xZnxj0o
InrKquhOTW1bdKNP1ZsyXV8vsEb+jyE520erCKvrpFKU/0X0X5boAQiJRfEgPeyl2H8V2oYbeznn
pnrPTWaVOQC76XVVP89KlzftfkY65G2oPqpl+wpOQmLHP8mCgVWVrd0B+qfH1wCuLBZ8gAYBsDl5
Abkgc7u1+jAJbAaR1k1IBV8j4qrnwpeJVSXqMu737otlrNpnMQy6m+O4GyYwlVlZLXENRQltIZMQ
i56+BKAmph2ittkHWqo/ahDME68Sz1E2JaikoI8xoe5o9L/5IPNVMkfM0WaeOioBXBQJ0FweLTYS
oeC+UE4qoFhF5+ohwkgJCXPbdRoGF4rk8C5N1fk5tKiamrWxNd9TOxew62/7byERAZtCkJsfg4f5
A5BLQQF7wXnBMfweP3ax5dwSvKczIDOCg3SkCFHMvqm00ea1ZfzLHCO/BkwqPVpvc0enG+Akz3AU
ro8RlAJ1W/xW+b0cYRogrfCRW353TI5DSZm7FzJ10Yl+o/JVLuGvX6lxpETBFb3BX9W3DSerSBAz
JcPj2Sk50y++oQ5wOpLl/ueqlGjQKVqh+YRmS3tHjC2hW1UE+vl7Nm/s/xrLTd+BkzIhR7Kq8CnL
8Aq4yYg21JCiDNTxhF99J62WUaVwPprREXFQp1cWzyA/AE6quN6DvmS7gRcBmpchmoOKI3vrnfMM
kqNn0wPfa2Gqb+3qHelruMezOCRcWJVMxrEv6e1ZRtLJluptgQ1eO5a3kdtxnSP8zBytSVdPVTQM
3Anc1F33Nm8WxpEV3W78cuxH4TZP6P3aBEJ2zG0AMg+og7I8SbYNv7BRBZP7gWFNzyy7f2DhlQwj
DLK2IJH3jZhEsL+n06CV7DNoKbOo1s7Phmbkn5Z2VKj6tStfQe/LBnd+hDTeG747XQSR4pIstNEI
YtFlemvQRR/pgzb82/od4h3tFTiw1EcODorRUounpy5BsIknMrUbvfcTpKxDSKvrAqNdA5zsag2p
bnt8bmtahP/+5bRTnefY5cdRkSs8wmDU+iQ65xTo5F3C6n/XaysEHP3BHWwQiQHqFwcc4IfQ4yeI
X6A6eOzfSWXZr4IgVURR2zG0WDtGfV18cr0L3/ODKDpBS4wmCkhqIq9LQbCC1VQ7yGK7IO8u5PrI
TWw6brUtEGuRUmkGRB69X+mnNIWdD5v4zmsrJof4BBYzX1SlKLMUC0Q3YDU6AlcA09zWBy/+RCvL
NIkEg7uWdZ7P6QCBTVg+CItse7+sKkzk5qZ0q8r6LtbpiNma5S9HwkxpPU0ZRpNbAH7FTyYbYGBQ
beMlNvAntR44oTRtasJI6S91lps3bpjG8aARf6XRmYJyLg+AWScztCWistxQu0YPCGg1o8jehiV9
2A2i9FBQ4v+vnl4VLCUVvu/vTJAlnjd+uDGjBoq9NFbmlPOZthI04osJ6rgYOeGTjQLMysD0L8Jb
+1QcGSlBd0lSGZr2ZbH0QeAPEvyNRls9F3f/DZM6y80Nf41jfVq64gc8G1BDuCr+v83XlyJLTj9N
XaXYk+PhC9w21Io6rQiNELn7XZBUH0bjgRyTtKg957Sy3PKlmyUbLAYnsqdnj5QzO1dLHu6qvtB0
CKd9crozLy4PBaGpDhTfBMuqfcBzSeFOYEsjHE1Utz76VTzXZRqHrE0dvJZqkM62nZ1AkN9XXFqR
y/b2JLtFSBhPN6RIfOOHpEx/as21oFz3ccmAyAogJgGvaRWkTZlt8AxCdVFSH+HXoYwqvOwXaVSG
vPhsrOMQBBjXnRbL1oUIXu2LwYcT0eFzTbtWOh/OI4AMm6kUcTNHT2gCuPDgbaOKEUVHaNNU8kPY
VL8Wd0Py0LnQgKXiMdSEkU7psC3MTz3QumScjgsTlpqHr/J5zA7BTU45qIRjmXQYvfTXEnt0j0Vw
J+4ktM1VFZi1PMAGMcBJhlaLAkh2qLTj8QUOhS9UGWW+PT5TXzjQqugcL6kuH2ByeC1Fm8rNneJp
8YBAFhRbFo/gtqWo90eH7im+6aVRqerIqB36LxujNolgVusYlVrtBpZpkO+VjRqx67oqCD1ci6GR
jd/pQXuWAj80MYc7lF9DGgg72ySusqjXba3yeaTIjYyZNQHf8UTzy+dHcuMEtSTv55jjXREqUDfV
uGj7MXr7B4Y/KdQZm2jtOn9RXG1Jlbv3uZ2sxs05qpN3zmCUbxk/KcuDgDmPgItIcOuI8zbNctPE
dZS6V4pUqOwFklbM5GmRE7kIOK5ks1JNwihoUn/CKrcD5fdv13v35PgVxqsFh6uucGdWW7UAmgZ+
Fz03A0ktXFNYoxNcPd56IDlsgNmaQ3sQvQvMas6c6bXPQdiJvf7jbIrjvfr5Udk84BHBajuTRGRt
WYn0OTRLR0hrkxbMkvfyNBcZEQyug3HSPSZc2fpCc+LlIviSmjrJ+fLSO1ifHpO60x+l6FNTXrXc
Ta5jliOfT5Mp9OmKz8zRwYcHaNVen2zMSDzKdzEAcUbsUnzfrYYJefgtWOVKB1YHTmH/MW40fRIl
S9n6woj2vIxSk5ugWaB/mM4ngFMSuj00NBO9MYBpsS/p/8Nm6OZF41REsnyqPqeiMQpBCouLpPx1
jaiyLau7dUyJimZ9L33bL5M73/cSuhv6zK09vkI8JhaIyOMJsUyDFQwN2BuxRlQ7gCcYpSTEHGNu
mMHiFVf+8X93810aS68bCwCJy09JGwqy2XaZn02bhyruIF6pKcuM08ipQ1Y0ufDceTnReYOT1gIO
Iy9thjxQHNx1Npd/OfGIBC3fEHXwwaCD5uxno2RqpaZMROdBOq72wy85UncsVE9QhWKfLMFa/Q8d
QPtauSfQXtLhe2v9OUWYDNh3RvhZ0SyIjHOJIrkSM4CIIUuidnNAdNlZdkAZtEZ0/lh8xZItmVAB
KaTw6aNx0YWXdSuSryuwmeEpIGAwhft3Dsmjt6zGQbNarQ2NjfRdKy0xipD/eWCUT4iplLAsIwan
+4+viWbgxICwH2xUNs0gjQKW28BmHiMm+Meo91gqYgZ/8IDPeSSXHA41vBI4BLOrvcDfMhfAmmDu
W8tafTr827gZonZN2KNP0y47L0wf3is2VQLdvl2TLs7FqzfmoBqnwjqm1uo1DZLEmoTEHSib/DQC
LghbdAnYq0l/11SX76+SQE3HnEIb/tU9H6HludYpHmtCwXBLH8KRDDAy0TMNw5ltqZO+XLzC6JlC
WctmfGDzI/qJrL1rImyWZar3hzWSP3KPGqQjWXFPzCDe07heR6M/wnGnX4D6gKQ4BKVQf0dQYOit
u9IpFMM5NxKfygLMOrxAGnxxizuiqDK3Ld7kowZ7dPOKT5IZ1Vb+0uqYKpTbAUIW0zAKsfhnrRx6
AtGdg1e/TowS/kp53GZuAFoEpOJQdSBnH+DJEgGqtyYTvbk1GJd3M61vApWEJTzWhreO+I3NqEj6
isvVuEkWFdHjc5Zr8Oae7oIiXjK0DRFXaDiM4AR1E7YVBeXui5EkOl24jh29hN9ajZ3bG8YPtovU
OHiWoH8snK5j9oule1B0tM88L/EF4waIGp7Asna1f/0ENH4eWABX6bJdKQJjkJu8BBTTjlV3t00r
tbLJY81xW5xnCcjDWzInSg6UnoxfJgJV6W/hcyUI/h6BQAzn2eaWV2QZvarvrzRedW831TbG7wIT
njt2BEuWsspDESsdqBRW/qInzLWsfBKnk7L0YYS/AuTWrg0OqEqOWocQQzIfLfFJD7JlGXQYKFDA
/+PV7KPN3GdLciF7AOsi1XVQfjVZ+p5WP5UCOdv4dmsoVzYWXbtS3fomjhb5sRhZkiVVesa3wmih
aNVPq3pt0M21ra88UuRe8AehJeC1Creu5SB7/O/fNx/4hloVMHSpEyLsjGQzPo7e0WWYu7r8pqlc
w4lyDfsLhbn8STh9EnfDmC3xh9NogA8Ida9PwyOaWEFucfb5rgpCgFE5CSLq7tQ87Geq3blyBuUG
4F6R8cWgHiY6PeQhPzB44gmxVkH9zp4KFskZaNyk6MJyapWQgIqo4tn+yU6JVgLF7Ug1PTE9f2pK
PjliFQscuZO4STl8xQgwX+kwII1OPE3qn3eb0DyZ9kvu/aH49nCLF0humE6fB4r6sQtoU7Q1o1Ap
FuIS7Y9BauqonENrTYK22r9nHr1n2aRJe1zaPGH2K+lowmNGQHUyM0rMiVg1SwYigi6v1RuZ8Wh7
uLYLyktypg+p1xh3n4NPqydI/Y9cTeH5mKaRC/58iArtYfjJK569hj58w1qGW8jMIL24BCS8myr9
IgSGeWzRrNJyskyNqSCAGTnQadXt8okrlL98V+IPCqN5MOd2e0G+hBgdNO2c+W9Rr+46xzHO3t2T
huKpHKBjxd8G5H1mBnLB62hub4EDxGVzQvcnwFohFf1+/69Hiv13TN97vzi9CBeKKNxBv9vrS4vB
wm73dUbJB6ikO0c2iJ45U3oMcC/gyw/8CxM371BpdVd/SaIkejN9IqI9YADbxTrIkqJBGMcvpPBx
WoSxkbWa6LOk/q6YDhpQ0o37+CAMvrJSpRX5vrTp4s6lIZ2VIXDd+YQUeEICLa5YydUWfLImn7bW
xbvHTZd/qo5/dELN/+TlFNjH+AuM4kWEMVqwlWQ3gUKXawX0rTghyltsDBAqpYI/LAQgfBHtIo5X
A4akWgrMG02xOzNcBaw5V3d95qphOWnxUpndoEx9dhP/TXVXEWGdE4hJpN10T+QBiIxKpk5HaLgg
cMJKuBV/eR94aHCk7T83S6q6EXArYYS2RNpwPECBy9HG46Prrqe9TJVClJpNq5leoEPo5kqZu1dz
Y84Uu+8dlORn7vl7K0KNgHf8DI76DCHYxSJHO/sd2vpB/cFQQTHrjSz1lL9LTEAmWCmMwxt61OLQ
lTPsCjvfjAelBf6loq3Ryvl+hp4zgUn9TN9SbzDM7P2Eeze95JXtIouBYoVGH337W/L7WrRbu5X6
zwNP2EZI/N5mbRgm3IaZUg2ev88OtKzY3vTBMOXvj+lf+5SrcEZQmiRcLX2PcSALhAiURbD8fxiW
qROTrWLAQ38Xrwuy+CBcwm5E/2ApeOFL/lO3fEa31wURra6zAJlOGMYNBoL847Urnba3gFygyUCV
cO+v1JPBBS/w5bZdPqEo05EbPigzxIWaYpSGf/QWM3J8nxxm9h8FvCfoI80RUDPwWrVdb6oPsE4R
Gxdw+aulwM0/GLhotKvZGbLCmNsDDE+VnD/i2mqjaG+yTFbdDZsoajkX3pgNpGPcwXh/4ycXz5hP
Yo4p9fuYIRYncYBGb0+PIfKm4c6lbpWiqorhljui/NWfnJmPk/vni0T0vBfMnrK8roRwI1GbIaow
3WC0yAnDiEHKoS4I5gIy/tbRSb77+DVmnGt+TIuHUtvk4dkcpKZRi4E4wl1AS4iOZAUgU4AUNtYx
94c4eD3qSOKpZ3TpmbDHZC6jRNhT4yTHofFJ06WO7lqI0C7jvNcQT6PH0/a4Qh1SEKS5mBH5Ful0
dBCgJdbXEUu/y9H0ca54x2KY09+6lzJDZx1efgoCWarJ9rfy+h6EP9Eib8n4UnHszIKiynz7J15r
ZugXd4uVYjkqOpVj2ZnmGuGRiL7myZCoIh1F8iMJ1ETHAf+ngslNvmftoJC1siYtOD/WhkwGQrbx
VK55mamdQW5+IfNFymvZkq+ETstjCDcLdIRHWfdSrzdDNBRqCoN9cD0ddXUrNALDJCtzFzDJcjRa
qf7uYYumBQBU+1+fKWQ7y2JYqwiLtvQVy9Mii87tomJyQDV4KwOxg0P6yKJ/mhRDt3w4p/oEBf21
qjvDdaWAqXmLPTBQJwiX/zak8V0mAdSaaYF6HdhM371pWmc8nhXg73p9eXS+CyqtTYRVmvxvgA39
EOd8s29+Teri6U7F708ZUXcSdZ+Jwq6mh4GC0HDgJkublz6FLKQ7jLbLPvZYhgaWVgLWjl9UAawb
paY09H7dr/+yZ24yGWuN9KUeTWhLnf2DOx7lGufaoCGB5DgSsBkso1a5AdWsDG3vJpaigqw6Dgl4
uyH9oDKHJ/EDhqKX3Uem98xpR6ti6+//q3jNjCUvQNwb2NIfXMJua+JTSAf+Qc2/YUdIPjUYqeN0
MGjoPmljPpSNSPKVl8kspgzRXCzJXIA7jAuW1/EL7P0YlZkp6xDrYRviLmoc0Ze9xY5yUFcRwTlV
GktNhMNq54CcPp2fDXhz4bnPHwqlJokXtPqLpEucmw4xDQj4j/l5gK0doHQ5Q4yEot4OQqvlKl6w
QIrBQJ5UWIJ8sT06kLA/cgpPWwSNrH6emiCRZA0VdaSs8TuOGmEUkly6yDKcysTbITXvcb3AMPpQ
6SRZ89cLrp2NtJRbBZ5D1iou/ztUECM8pITGOE8pLsmT/mfyngSYR/LV9snP2qoaUwaLR8A/mPHB
IhwZ/1EsUpxQDquQ3MkEo1ZD2X/51NJVmmwe31pZYWZOBa4UF1frX6hS2QzVh4hTrbWpTqYED1da
/TX8H+t+pMxAlVTtpyOdX/nVPpfNH5UTP3G2gj3L23BaPdYyjnsjpDJFkxsY0j8t3BlxEr8qwzPJ
fPUQ/HzujHdFuzKx3kXu3KPhtQhteAlOWU2NpFrjYh6+96PZz2yEw9rD4zIqE7FiXdM0L2ny/S0B
gtMi5Fx+SCpx/H+XwtMITUCRPe0p1OxVd9Lk5oFVGsP+WkDRzdywrH8Z9Ha+sonHkfrSrBwCCO9y
SxWthIeLEzyDya3YzWBScCtc4eWKWQAm9YgM81LmSHjWiq9os9HS0hfuLQUW42AEjEZZpO9YUKi3
4e7kMlBDXg0eK0tf7hO6WThk4QYvHyEfw+bUaVrJ1cSr1L/YhMCgGbShOq8cBgjM84dhzBN028y7
qZhK8gcHc415ul/UQcZ5TepxWEH2H+EZ13el4wjfzgh+5jeEorDHneuZf+KTo1VSaWGUJjhDDHHX
piPdKxx7JDNMy4t/E3EV3pvVdfOxNhOtVEdzs+zSprHifM2Y+jxCwsM5jW2dD4T+YjDNDjmfi5w8
Clo6Q2kcWKk0QRnzTab+UG91xZyeAyie2Yto3Q1GS1pFxKB87n3LU9nWJJ7gaLgvvRJQ60CNRrXq
1L6Z9+gMvHbZyThUImu12cTtDmxjsQU14lUtVMzRDe3CD4h0gqk2DrzUOctgzbslbf9LPblne0oD
a+gT+SLZq20hRo4ClHEvfwQqkC+PguKIhg0PtuNHxqk76dhAVcFqTPK2tHa5ad/XTQQvXSzWiSW3
0Ea/J1kNzVHfPnC5mD55DTKV7IhDH2vbSEYLZNtXmJxvbuc6GH9HPIPnVe3on6XFcr9It5ahdeds
5GFgbEvxQZ5sg/2wbDyPtO5SBPocZDLITDjoxWyJIGEGviPY3gpWlBVgf312Q9JYBPM/DfC5QrqJ
Py6Bpbys+p6aSLpAPrdrEHELY+FZ78oGnTnG2tEW/Qep8lAD5QUsdskrAUZF1y6h5wEUBgiIjoK7
ibZi4dkLU/1Zn0lrHy6hwLrIvYiKLOJMpn/LIW/hWIE2BAOxpAwb8NcbBB990pDHc+/t5LnMUrZ3
wVWvbbX8xLZAo2cvUA4yCddFqTu5YgdSE+pIcGMiAxLV/gattv/co/YkPawxjwMM676Mu+uzHG74
sxxONKzo/AAUMFlPw08l3HOwPaH3wKJG0sHqR3vnbHYNkl48Vv71QWg9Ks4owQS/L3ciiBS9+NC6
jSn3PYw/ZKoFCHJBkAWvItm2/FE9swhz4K7fWL5KG4xkA5gjlVsEOv/P8Bh/GrQBfPVjIrQDJ+E6
frL1P6u7kD2u/RTogQuFjZouz4SwsJzKZeHX/zChy0puxGowLYGfHnT5aHFL+o6hjEPh7hvRh7My
WzlQMHNLklLzu+AQ62YoP1qPQZqTDsKSujvIvUP1IfMf8wyxE8bNnDw58Rfq0I/A9xJtc/Gcao2k
mshvUP3Zk3ttcHJmWrC1Bt0ETzZ7p+Zqt2WzANJNRmtYsfFmTYiUS5tETOojqSJE+fbaf2Kh2MxB
03ACD7fmTpNDxWUz4IHAwXRdP4kFE+p/auur9eEur6PMpPvOU3fy2ZeyQONYYnz2//qzFOJs6GYo
hrJ4caajvO+RiQtFm1H6t8quaV7+OPQY67NIg+xydHDSc7B1ZHjppH2YKnAiyoKJrfsjJqkMV6sq
3LJnrzt9MGZwQOp2UekEgnFVsdsYFXzdLxa8H8XO43o5KBnqpVE0byR7GU32eELcYkr9SSCjJj76
F+PQ1yt9JLlFk3Di6Wtk9T5kblly6YL53XvFPzOq3G0jlwH3dJ6wpb8Kf4xalkIyPWvoR5USaG5f
/4Svhrs24Zfg5DGNsfqRai/mWcL1ICKvbfUboDQcszrHWjPtit2Uhvusm+lQPz7h4tY1nlU6SAjc
wsB/+I3zTjGTUOXZppjzGJWyiZ8hzvUsPvPU28S4tPa67slJv2rXf6dmFe9fz52XOV1wASI4GLA2
cRkoo6J+znVf4haZ2cNERryRMMz62nTfnjj1hwpt4zKsVvOIFqsLFEacY+A+c74sr9jk+KQ2p1fC
9HCZrbC3XgTCQkiTY9SSp0qtMemx0fLArd372YgGEeu/pnKMDGL/sXTLl8Ja9nv9f937KAs5Dhda
0B2spzxYBulaFPBRkZydJ6iSQofdt2bwjwDxg7QDJS9McjquYlpBq4ktTHbARcsx6xpHLEfKsq1Z
YZWsXnGLYUHFrWgYj3Z0R9ihbe9vW6XGbhUTqz25EloUMYsXMmE1D/49+LZmZsh8yJ28ZvyicgyA
dOnQfGN9UAVFzJAwF7YmsxgJpNteFkc1ahONutl0Js/Q2OB+AiorBVH699DFwKYZ1wNjDIzG5sND
jkkNZouEhxJ8MpFP6rn4569VK6D05em6kK59hXyY021jvRNuM5XI3N4LAWtxhXjENc9SViqOIufC
M7NqoIqSWjy3nImwXcMRbenfdMTpoVR/38BSBD91piJUo7beVGhc3eFGiDOHhGOmq8OkJGGuJpjY
yXKl+lXSSj7DJbiBhrdirNqYNmz90a9Yv+6nECh3kz2gHa13sKNuys+1K9melaq8ntJZIQcZ59sU
uVbxEa0LxtEvcWVlK8wOXaSfMynLnMqX5ydMAgN68bim/7UmOmmANNwD5Y5TfCa8CfdOt8fxTPqk
h3IX07DbqjOdj6lvEFvqZij6knIxL/bDGg7YEPnSak3Eg40cRCnzIh4OXpNzuIHkSAL0h3AxESLb
00w41i+4/6+6l7HDPQjiKuCSk6PwLjo9QAokvdujWLmvH+G78OvGlhh1Omr+gwrVr2IW18nUZe4z
niJzUV1TOoYt5JcaLjWoNMzmb37zAS94jzPs2J/Tfs0RgfmTAFd1vP1R0RcCesUfFUksX6QTZecZ
j8L2tFWd0yEKYVIllWRM4F6jVUnPmjgyKHJXpz/AMPQ48GO1r5+kipLsz73aRNOGykYpmpwDkY7M
gAAG0dLgeWdCse18ramRxZ6mgHygDlpFJWwSjeHBcsNq9gHlnkzpa5GJrFavXuW/zeNMCr8V+UMi
s+019EgVKCNyIL4Qam1NtN/FSbKDV2eMMyz1REY/8ai5jwTJT6iaultnssLfqB294NfOt1/Q57Rt
nhbb9d184zqfSifiqTl6R1k0hqPPvFUFcWfpA3YoOFXillMOT/ny5pdvV76YQSF04N0RCpph8+Cn
E73ZDFuEoJL2/sttNqblzdwhlnM+LnIlqbPTJyBD6InHiL95H21BpuYTVfgbFjxCDoS/I48p9ed8
+kWEQFnAldN+ES7dZIfKLYhZPo2WKATDht85hOe2KzIuTrZf9WhHbjUzroxD5nqGTyRhcbBhZkUb
EvlU2aCBFl3Kxfz1FGwNA4cH8IFV0jw4fAdhN8bmW2RsWp+o95tF7xhyc5kM4Os63Mb7i7hfodgU
y60g2LKisTOX1wVg0FaHVaYo8UPFIIoTkp+NINoa/mVQs3OF7wSTWMllOhuIhUDQ1mLH+uYjXAvy
lpFbdPOrBBCzUYqlwKLJ/K8XwusAcSEFjKNI/Fbhq8om/TEmVApilMuF842L/ya6OsUeW2drZLsU
azBlnqH8ixB3Cp9dbXOujIsnUN1b3VojttppJQs4S3KzkxIffr08ZC5qoKzK4GLOc0lY8wb52n0N
vET9EFsXvMlhTNFAMPbp4D6wDyzeR5WEHeB4wcvQL7k+B5ruB8Q0F4KtYURfI3IQrfjKiUZprtcJ
RzNt4U1SOM4pJpOkISZixSGzu806pfdP2NaXhQ6FcdsiqwYC0bGtUQzG6QFZcNnCuTfXH25heIJt
LAm8MuRJKQRxsW28B3tUhA4O7OxvJRWXsf+Pz+xiRHS/zgWQK1rV5yR4bBFyiQLLU5Os10FB9vbG
lffR7Oer3cREdpRFevp6Ge261ghNZgM4e+h/ewkUkpt/GLc5En4dFFepaFu7m3RUOZZlCIW3Iz9b
BVNoBZh9+Jl7C8FvAy8F2o/YAWsA2WfX9tiBz0XpWiQNGV0QWGbH6kkORNOiVmtKl3bbIjguTEU9
+dxJAzDCEVN7FqS+CgqcwEpX020s1luX8JbzFRqrbfkt8ElhuvqkD5AxB5FhZODlCFeTeUBhhXGV
f8AS4VMg8ocyPetMm1vtogb/fTWFbbE4qDVM+M6BxByia05XMjFaBqwPumKnj2MTHFOzVOkoEbdm
vUYQQ8w/aRTT7ZqD18PQhWMh4AOgxo8XI3hLfz333QRgH+6xFVTvMpQ6+kCQvwBc32krvU9/qPnk
6xD47/ycPlH5BoG7eLKmvI6JCyydVeI1WmZh1r1JkkFxc6rFwq+kZ1MVtVFVpD+DBYOto43W1f7u
gY4MG+F3CaOOycK2ize9YlbEigyeeapIengb2l4g0UiPskWxzdS36V3BnC+XU2Nu9/xcQ+cVkYf3
rmaAsV6HdjKR2leJSnUewYaIVk/i5K63f1lCHVCMX9e2307XuIAk/XpDTB8GXFs3Hbi5K/H6+zMz
6StZpf4c9DVeeA8bFNZ2sQVmp17TcEfT5XpWUZZSy9rYhulMoUAh/sB4hulxXbNCmPjGySNhXfLi
fIMdIRoH2K/bF0lCzmXcrSCqNp5uaYFTpME3N+8VO+j2db8evSVyU0Ywl46EjMdpQllShy7Y0/DR
FR4Wz931yGewWARRfbT6rnQ+NyXlreE67dx/0pmSKqlYcIO124GR4TxcXa6718/ZCQEpNFC6BKwy
4KnK441wWIjEK3S7i/b3EsgP0+JYAVa3ySGOJVopIUsdrJGAfWSEffaJlkPgMwA/K9cgRoDeHDmd
hXldgF4WA3s9MRRnHWX0FlxcjoNqd8GwLJ5BfWbcKWsG5Lq+PdiK4JUHdjX7En6BV2SKcS1RoMBo
XoMsmuoO/NaZadXzpz2F6ksbCi3NgqXZiNNxrlOgkRSHphynFcsLneJaIwx2Hk12VOivUaxM+m2f
pmL8hV0a9PRpPmptxf5h5ZsZ1yBViVgP3EzCXDYpA5Dw0a2BQUYDtNvgRtfkXC5LbbtKh9dLfdmz
Y90tS0ogAS8Y8oX1aYQ=
`protect end_protected
